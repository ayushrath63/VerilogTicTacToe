module grid_rom(
//inputs
clk, addr, 
//outputs
data);

(* rom_style = "block" *)

input wire clk;
input wire [15:0] addr;
output reg [7:0] data = 0;

reg [15:0] addr_reg;

always @ (posedge clk)
	addr_reg <= addr;

always @ (*)
begin
	case(addr)
		16'b0000000001001110: data <= 8'b11111111;
		16'b0000000001001111: data <= 8'b11111111;
		16'b0000000001010000: data <= 8'b11111111;
		16'b0000000001010001: data <= 8'b11111111;
		16'b0000000010011110: data <= 8'b11111111;
		16'b0000000010011111: data <= 8'b11111111;
		16'b0000000010100000: data <= 8'b11111111;
		16'b0000000010100001: data <= 8'b11111111;
		16'b0000000100111110: data <= 8'b11111111;
		16'b0000000100111111: data <= 8'b11111111;
		16'b0000000101000000: data <= 8'b11111111;
		16'b0000000101000001: data <= 8'b11111111;
		16'b0000000110001110: data <= 8'b11111111;
		16'b0000000110001111: data <= 8'b11111111;
		16'b0000000110010000: data <= 8'b11111111;
		16'b0000000110010001: data <= 8'b11111111;
		16'b0000001000101110: data <= 8'b11111111;
		16'b0000001000101111: data <= 8'b11111111;
		16'b0000001000110000: data <= 8'b11111111;
		16'b0000001000110001: data <= 8'b11111111;
		16'b0000001001111110: data <= 8'b11111111;
		16'b0000001001111111: data <= 8'b11111111;
		16'b0000001010000000: data <= 8'b11111111;
		16'b0000001010000001: data <= 8'b11111111;
		16'b0000001100011110: data <= 8'b11111111;
		16'b0000001100011111: data <= 8'b11111111;
		16'b0000001100100000: data <= 8'b11111111;
		16'b0000001100100001: data <= 8'b11111111;
		16'b0000001101101110: data <= 8'b11111111;
		16'b0000001101101111: data <= 8'b11111111;
		16'b0000001101110000: data <= 8'b11111111;
		16'b0000001101110001: data <= 8'b11111111;
		16'b0000010000001110: data <= 8'b11111111;
		16'b0000010000001111: data <= 8'b11111111;
		16'b0000010000010000: data <= 8'b11111111;
		16'b0000010000010001: data <= 8'b11111111;
		16'b0000010001011110: data <= 8'b11111111;
		16'b0000010001011111: data <= 8'b11111111;
		16'b0000010001100000: data <= 8'b11111111;
		16'b0000010001100001: data <= 8'b11111111;
		16'b0000010011111110: data <= 8'b11111111;
		16'b0000010011111111: data <= 8'b11111111;
		16'b0000010100000000: data <= 8'b11111111;
		16'b0000010100000001: data <= 8'b11111111;
		16'b0000010101001110: data <= 8'b11111111;
		16'b0000010101001111: data <= 8'b11111111;
		16'b0000010101010000: data <= 8'b11111111;
		16'b0000010101010001: data <= 8'b11111111;
		16'b0000010111101110: data <= 8'b11111111;
		16'b0000010111101111: data <= 8'b11111111;
		16'b0000010111110000: data <= 8'b11111111;
		16'b0000010111110001: data <= 8'b11111111;
		16'b0000011000111110: data <= 8'b11111111;
		16'b0000011000111111: data <= 8'b11111111;
		16'b0000011001000000: data <= 8'b11111111;
		16'b0000011001000001: data <= 8'b11111111;
		16'b0000011011011110: data <= 8'b11111111;
		16'b0000011011011111: data <= 8'b11111111;
		16'b0000011011100000: data <= 8'b11111111;
		16'b0000011011100001: data <= 8'b11111111;
		16'b0000011100101110: data <= 8'b11111111;
		16'b0000011100101111: data <= 8'b11111111;
		16'b0000011100110000: data <= 8'b11111111;
		16'b0000011100110001: data <= 8'b11111111;
		16'b0000011111001110: data <= 8'b11111111;
		16'b0000011111001111: data <= 8'b11111111;
		16'b0000011111010000: data <= 8'b11111111;
		16'b0000011111010001: data <= 8'b11111111;
		16'b0000100000011110: data <= 8'b11111111;
		16'b0000100000011111: data <= 8'b11111111;
		16'b0000100000100000: data <= 8'b11111111;
		16'b0000100000100001: data <= 8'b11111111;
		16'b0000100010111110: data <= 8'b11111111;
		16'b0000100010111111: data <= 8'b11111111;
		16'b0000100011000000: data <= 8'b11111111;
		16'b0000100011000001: data <= 8'b11111111;
		16'b0000100100001110: data <= 8'b11111111;
		16'b0000100100001111: data <= 8'b11111111;
		16'b0000100100010000: data <= 8'b11111111;
		16'b0000100100010001: data <= 8'b11111111;
		16'b0000100110101110: data <= 8'b11111111;
		16'b0000100110101111: data <= 8'b11111111;
		16'b0000100110110000: data <= 8'b11111111;
		16'b0000100110110001: data <= 8'b11111111;
		16'b0000100111111110: data <= 8'b11111111;
		16'b0000100111111111: data <= 8'b11111111;
		16'b0000101000000000: data <= 8'b11111111;
		16'b0000101000000001: data <= 8'b11111111;
		16'b0000101010011110: data <= 8'b11111111;
		16'b0000101010011111: data <= 8'b11111111;
		16'b0000101010100000: data <= 8'b11111111;
		16'b0000101010100001: data <= 8'b11111111;
		16'b0000101011101110: data <= 8'b11111111;
		16'b0000101011101111: data <= 8'b11111111;
		16'b0000101011110000: data <= 8'b11111111;
		16'b0000101011110001: data <= 8'b11111111;
		16'b0000101110001110: data <= 8'b11111111;
		16'b0000101110001111: data <= 8'b11111111;
		16'b0000101110010000: data <= 8'b11111111;
		16'b0000101110010001: data <= 8'b11111111;
		16'b0000101111011110: data <= 8'b11111111;
		16'b0000101111011111: data <= 8'b11111111;
		16'b0000101111100000: data <= 8'b11111111;
		16'b0000101111100001: data <= 8'b11111111;
		16'b0000110001111110: data <= 8'b11111111;
		16'b0000110001111111: data <= 8'b11111111;
		16'b0000110010000000: data <= 8'b11111111;
		16'b0000110010000001: data <= 8'b11111111;
		16'b0000110011001110: data <= 8'b11111111;
		16'b0000110011001111: data <= 8'b11111111;
		16'b0000110011010000: data <= 8'b11111111;
		16'b0000110011010001: data <= 8'b11111111;
		16'b0000110101101110: data <= 8'b11111111;
		16'b0000110101101111: data <= 8'b11111111;
		16'b0000110101110000: data <= 8'b11111111;
		16'b0000110101110001: data <= 8'b11111111;
		16'b0000110110111110: data <= 8'b11111111;
		16'b0000110110111111: data <= 8'b11111111;
		16'b0000110111000000: data <= 8'b11111111;
		16'b0000110111000001: data <= 8'b11111111;
		16'b0000111001011110: data <= 8'b11111111;
		16'b0000111001011111: data <= 8'b11111111;
		16'b0000111001100000: data <= 8'b11111111;
		16'b0000111001100001: data <= 8'b11111111;
		16'b0000111010101110: data <= 8'b11111111;
		16'b0000111010101111: data <= 8'b11111111;
		16'b0000111010110000: data <= 8'b11111111;
		16'b0000111010110001: data <= 8'b11111111;
		16'b0000111101001110: data <= 8'b11111111;
		16'b0000111101001111: data <= 8'b11111111;
		16'b0000111101010000: data <= 8'b11111111;
		16'b0000111101010001: data <= 8'b11111111;
		16'b0000111110011110: data <= 8'b11111111;
		16'b0000111110011111: data <= 8'b11111111;
		16'b0000111110100000: data <= 8'b11111111;
		16'b0000111110100001: data <= 8'b11111111;
		16'b0001000000111110: data <= 8'b11111111;
		16'b0001000000111111: data <= 8'b11111111;
		16'b0001000001000000: data <= 8'b11111111;
		16'b0001000001000001: data <= 8'b11111111;
		16'b0001000010001110: data <= 8'b11111111;
		16'b0001000010001111: data <= 8'b11111111;
		16'b0001000010010000: data <= 8'b11111111;
		16'b0001000010010001: data <= 8'b11111111;
		16'b0001000100101110: data <= 8'b11111111;
		16'b0001000100101111: data <= 8'b11111111;
		16'b0001000100110000: data <= 8'b11111111;
		16'b0001000100110001: data <= 8'b11111111;
		16'b0001000101111110: data <= 8'b11111111;
		16'b0001000101111111: data <= 8'b11111111;
		16'b0001000110000000: data <= 8'b11111111;
		16'b0001000110000001: data <= 8'b11111111;
		16'b0001001000011110: data <= 8'b11111111;
		16'b0001001000011111: data <= 8'b11111111;
		16'b0001001000100000: data <= 8'b11111111;
		16'b0001001000100001: data <= 8'b11111111;
		16'b0001001001101110: data <= 8'b11111111;
		16'b0001001001101111: data <= 8'b11111111;
		16'b0001001001110000: data <= 8'b11111111;
		16'b0001001001110001: data <= 8'b11111111;
		16'b0001001100001110: data <= 8'b11111111;
		16'b0001001100001111: data <= 8'b11111111;
		16'b0001001100010000: data <= 8'b11111111;
		16'b0001001100010001: data <= 8'b11111111;
		16'b0001001101011110: data <= 8'b11111111;
		16'b0001001101011111: data <= 8'b11111111;
		16'b0001001101100000: data <= 8'b11111111;
		16'b0001001101100001: data <= 8'b11111111;
		16'b0001001111111110: data <= 8'b11111111;
		16'b0001001111111111: data <= 8'b11111111;
		16'b0001010000000000: data <= 8'b11111111;
		16'b0001010000000001: data <= 8'b11111111;
		16'b0001010001001110: data <= 8'b11111111;
		16'b0001010001001111: data <= 8'b11111111;
		16'b0001010001010000: data <= 8'b11111111;
		16'b0001010001010001: data <= 8'b11111111;
		16'b0001010011101110: data <= 8'b11111111;
		16'b0001010011101111: data <= 8'b11111111;
		16'b0001010011110000: data <= 8'b11111111;
		16'b0001010011110001: data <= 8'b11111111;
		16'b0001010100111110: data <= 8'b11111111;
		16'b0001010100111111: data <= 8'b11111111;
		16'b0001010101000000: data <= 8'b11111111;
		16'b0001010101000001: data <= 8'b11111111;
		16'b0001010111011110: data <= 8'b11111111;
		16'b0001010111011111: data <= 8'b11111111;
		16'b0001010111100000: data <= 8'b11111111;
		16'b0001010111100001: data <= 8'b11111111;
		16'b0001011000101110: data <= 8'b11111111;
		16'b0001011000101111: data <= 8'b11111111;
		16'b0001011000110000: data <= 8'b11111111;
		16'b0001011000110001: data <= 8'b11111111;
		16'b0001011011001110: data <= 8'b11111111;
		16'b0001011011001111: data <= 8'b11111111;
		16'b0001011011010000: data <= 8'b11111111;
		16'b0001011011010001: data <= 8'b11111111;
		16'b0001011100011110: data <= 8'b11111111;
		16'b0001011100011111: data <= 8'b11111111;
		16'b0001011100100000: data <= 8'b11111111;
		16'b0001011100100001: data <= 8'b11111111;
		16'b0001011110111110: data <= 8'b11111111;
		16'b0001011110111111: data <= 8'b11111111;
		16'b0001011111000000: data <= 8'b11111111;
		16'b0001011111000001: data <= 8'b11111111;
		16'b0001100000001110: data <= 8'b11111111;
		16'b0001100000001111: data <= 8'b11111111;
		16'b0001100000010000: data <= 8'b11111111;
		16'b0001100000010001: data <= 8'b11111111;
		16'b0001100010101110: data <= 8'b11111111;
		16'b0001100010101111: data <= 8'b11111111;
		16'b0001100010110000: data <= 8'b11111111;
		16'b0001100010110001: data <= 8'b11111111;
		16'b0001100011111110: data <= 8'b11111111;
		16'b0001100011111111: data <= 8'b11111111;
		16'b0001100100000000: data <= 8'b11111111;
		16'b0001100100000001: data <= 8'b11111111;
		16'b0001100110011110: data <= 8'b11111111;
		16'b0001100110011111: data <= 8'b11111111;
		16'b0001100110100000: data <= 8'b11111111;
		16'b0001100110100001: data <= 8'b11111111;
		16'b0001100111101110: data <= 8'b11111111;
		16'b0001100111101111: data <= 8'b11111111;
		16'b0001100111110000: data <= 8'b11111111;
		16'b0001100111110001: data <= 8'b11111111;
		16'b0001101010001110: data <= 8'b11111111;
		16'b0001101010001111: data <= 8'b11111111;
		16'b0001101010010000: data <= 8'b11111111;
		16'b0001101010010001: data <= 8'b11111111;
		16'b0001101011011110: data <= 8'b11111111;
		16'b0001101011011111: data <= 8'b11111111;
		16'b0001101011100000: data <= 8'b11111111;
		16'b0001101011100001: data <= 8'b11111111;
		16'b0001101101111110: data <= 8'b11111111;
		16'b0001101101111111: data <= 8'b11111111;
		16'b0001101110000000: data <= 8'b11111111;
		16'b0001101110000001: data <= 8'b11111111;
		16'b0001101111001110: data <= 8'b11111111;
		16'b0001101111001111: data <= 8'b11111111;
		16'b0001101111010000: data <= 8'b11111111;
		16'b0001101111010001: data <= 8'b11111111;
		16'b0001110001101110: data <= 8'b11111111;
		16'b0001110001101111: data <= 8'b11111111;
		16'b0001110001110000: data <= 8'b11111111;
		16'b0001110001110001: data <= 8'b11111111;
		16'b0001110010111110: data <= 8'b11111111;
		16'b0001110010111111: data <= 8'b11111111;
		16'b0001110011000000: data <= 8'b11111111;
		16'b0001110011000001: data <= 8'b11111111;
		16'b0001110101011110: data <= 8'b11111111;
		16'b0001110101011111: data <= 8'b11111111;
		16'b0001110101100000: data <= 8'b11111111;
		16'b0001110101100001: data <= 8'b11111111;
		16'b0001110110101110: data <= 8'b11111111;
		16'b0001110110101111: data <= 8'b11111111;
		16'b0001110110110000: data <= 8'b11111111;
		16'b0001110110110001: data <= 8'b11111111;
		16'b0001111001001110: data <= 8'b11111111;
		16'b0001111001001111: data <= 8'b11111111;
		16'b0001111001010000: data <= 8'b11111111;
		16'b0001111001010001: data <= 8'b11111111;
		16'b0001111010011110: data <= 8'b11111111;
		16'b0001111010011111: data <= 8'b11111111;
		16'b0001111010100000: data <= 8'b11111111;
		16'b0001111010100001: data <= 8'b11111111;
		16'b0001111100111110: data <= 8'b11111111;
		16'b0001111100111111: data <= 8'b11111111;
		16'b0001111101000000: data <= 8'b11111111;
		16'b0001111101000001: data <= 8'b11111111;
		16'b0001111110001110: data <= 8'b11111111;
		16'b0001111110001111: data <= 8'b11111111;
		16'b0001111110010000: data <= 8'b11111111;
		16'b0001111110010001: data <= 8'b11111111;
		16'b0010000000101110: data <= 8'b11111111;
		16'b0010000000101111: data <= 8'b11111111;
		16'b0010000000110000: data <= 8'b11111111;
		16'b0010000000110001: data <= 8'b11111111;
		16'b0010000001111110: data <= 8'b11111111;
		16'b0010000001111111: data <= 8'b11111111;
		16'b0010000010000000: data <= 8'b11111111;
		16'b0010000010000001: data <= 8'b11111111;
		16'b0010000100011110: data <= 8'b11111111;
		16'b0010000100011111: data <= 8'b11111111;
		16'b0010000100100000: data <= 8'b11111111;
		16'b0010000100100001: data <= 8'b11111111;
		16'b0010000101101110: data <= 8'b11111111;
		16'b0010000101101111: data <= 8'b11111111;
		16'b0010000101110000: data <= 8'b11111111;
		16'b0010000101110001: data <= 8'b11111111;
		16'b0010001000001110: data <= 8'b11111111;
		16'b0010001000001111: data <= 8'b11111111;
		16'b0010001000010000: data <= 8'b11111111;
		16'b0010001000010001: data <= 8'b11111111;
		16'b0010001001011110: data <= 8'b11111111;
		16'b0010001001011111: data <= 8'b11111111;
		16'b0010001001100000: data <= 8'b11111111;
		16'b0010001001100001: data <= 8'b11111111;
		16'b0010001011111110: data <= 8'b11111111;
		16'b0010001011111111: data <= 8'b11111111;
		16'b0010001100000000: data <= 8'b11111111;
		16'b0010001100000001: data <= 8'b11111111;
		16'b0010001101001110: data <= 8'b11111111;
		16'b0010001101001111: data <= 8'b11111111;
		16'b0010001101010000: data <= 8'b11111111;
		16'b0010001101010001: data <= 8'b11111111;
		16'b0010001111101110: data <= 8'b11111111;
		16'b0010001111101111: data <= 8'b11111111;
		16'b0010001111110000: data <= 8'b11111111;
		16'b0010001111110001: data <= 8'b11111111;
		16'b0010010000111110: data <= 8'b11111111;
		16'b0010010000111111: data <= 8'b11111111;
		16'b0010010001000000: data <= 8'b11111111;
		16'b0010010001000001: data <= 8'b11111111;
		16'b0010010011011110: data <= 8'b11111111;
		16'b0010010011011111: data <= 8'b11111111;
		16'b0010010011100000: data <= 8'b11111111;
		16'b0010010011100001: data <= 8'b11111111;
		16'b0010010100101110: data <= 8'b11111111;
		16'b0010010100101111: data <= 8'b11111111;
		16'b0010010100110000: data <= 8'b11111111;
		16'b0010010100110001: data <= 8'b11111111;
		16'b0010010111001110: data <= 8'b11111111;
		16'b0010010111001111: data <= 8'b11111111;
		16'b0010010111010000: data <= 8'b11111111;
		16'b0010010111010001: data <= 8'b11111111;
		16'b0010011000011110: data <= 8'b11111111;
		16'b0010011000011111: data <= 8'b11111111;
		16'b0010011000100000: data <= 8'b11111111;
		16'b0010011000100001: data <= 8'b11111111;
		16'b0010011010111110: data <= 8'b11111111;
		16'b0010011010111111: data <= 8'b11111111;
		16'b0010011011000000: data <= 8'b11111111;
		16'b0010011011000001: data <= 8'b11111111;
		16'b0010011100001110: data <= 8'b11111111;
		16'b0010011100001111: data <= 8'b11111111;
		16'b0010011100010000: data <= 8'b11111111;
		16'b0010011100010001: data <= 8'b11111111;
		16'b0010011110101110: data <= 8'b11111111;
		16'b0010011110101111: data <= 8'b11111111;
		16'b0010011110110000: data <= 8'b11111111;
		16'b0010011110110001: data <= 8'b11111111;
		16'b0010011111111110: data <= 8'b11111111;
		16'b0010011111111111: data <= 8'b11111111;
		16'b0010100000000000: data <= 8'b11111111;
		16'b0010100000000001: data <= 8'b11111111;
		16'b0010100010011110: data <= 8'b11111111;
		16'b0010100010011111: data <= 8'b11111111;
		16'b0010100010100000: data <= 8'b11111111;
		16'b0010100010100001: data <= 8'b11111111;
		16'b0010100011101110: data <= 8'b11111111;
		16'b0010100011101111: data <= 8'b11111111;
		16'b0010100011110000: data <= 8'b11111111;
		16'b0010100011110001: data <= 8'b11111111;
		16'b0010100110001110: data <= 8'b11111111;
		16'b0010100110001111: data <= 8'b11111111;
		16'b0010100110010000: data <= 8'b11111111;
		16'b0010100110010001: data <= 8'b11111111;
		16'b0010100111011110: data <= 8'b11111111;
		16'b0010100111011111: data <= 8'b11111111;
		16'b0010100111100000: data <= 8'b11111111;
		16'b0010100111100001: data <= 8'b11111111;
		16'b0010101001111110: data <= 8'b11111111;
		16'b0010101001111111: data <= 8'b11111111;
		16'b0010101010000000: data <= 8'b11111111;
		16'b0010101010000001: data <= 8'b11111111;
		16'b0010101011001110: data <= 8'b11111111;
		16'b0010101011001111: data <= 8'b11111111;
		16'b0010101011010000: data <= 8'b11111111;
		16'b0010101011010001: data <= 8'b11111111;
		16'b0010101101101110: data <= 8'b11111111;
		16'b0010101101101111: data <= 8'b11111111;
		16'b0010101101110000: data <= 8'b11111111;
		16'b0010101101110001: data <= 8'b11111111;
		16'b0010101110111110: data <= 8'b11111111;
		16'b0010101110111111: data <= 8'b11111111;
		16'b0010101111000000: data <= 8'b11111111;
		16'b0010101111000001: data <= 8'b11111111;
		16'b0010110001011110: data <= 8'b11111111;
		16'b0010110001011111: data <= 8'b11111111;
		16'b0010110001100000: data <= 8'b11111111;
		16'b0010110001100001: data <= 8'b11111111;
		16'b0010110010101110: data <= 8'b11111111;
		16'b0010110010101111: data <= 8'b11111111;
		16'b0010110010110000: data <= 8'b11111111;
		16'b0010110010110001: data <= 8'b11111111;
		16'b0010110101001110: data <= 8'b11111111;
		16'b0010110101001111: data <= 8'b11111111;
		16'b0010110101010000: data <= 8'b11111111;
		16'b0010110101010001: data <= 8'b11111111;
		16'b0010110110011110: data <= 8'b11111111;
		16'b0010110110011111: data <= 8'b11111111;
		16'b0010110110100000: data <= 8'b11111111;
		16'b0010110110100001: data <= 8'b11111111;
		16'b0010111000111110: data <= 8'b11111111;
		16'b0010111000111111: data <= 8'b11111111;
		16'b0010111001000000: data <= 8'b11111111;
		16'b0010111001000001: data <= 8'b11111111;
		16'b0010111010001110: data <= 8'b11111111;
		16'b0010111010001111: data <= 8'b11111111;
		16'b0010111010010000: data <= 8'b11111111;
		16'b0010111010010001: data <= 8'b11111111;
		16'b0010111100101110: data <= 8'b11111111;
		16'b0010111100101111: data <= 8'b11111111;
		16'b0010111100110000: data <= 8'b11111111;
		16'b0010111100110001: data <= 8'b11111111;
		16'b0010111101111110: data <= 8'b11111111;
		16'b0010111101111111: data <= 8'b11111111;
		16'b0010111110000000: data <= 8'b11111111;
		16'b0010111110000001: data <= 8'b11111111;
		16'b0011000000011110: data <= 8'b11111111;
		16'b0011000000011111: data <= 8'b11111111;
		16'b0011000000100000: data <= 8'b11111111;
		16'b0011000000100001: data <= 8'b11111111;
		16'b0011000001101110: data <= 8'b11111111;
		16'b0011000001101111: data <= 8'b11111111;
		16'b0011000001110000: data <= 8'b11111111;
		16'b0011000001110001: data <= 8'b11111111;
		16'b0011000100001110: data <= 8'b11111111;
		16'b0011000100001111: data <= 8'b11111111;
		16'b0011000100010000: data <= 8'b11111111;
		16'b0011000100010001: data <= 8'b11111111;
		16'b0011000101011110: data <= 8'b11111111;
		16'b0011000101011111: data <= 8'b11111111;
		16'b0011000101100000: data <= 8'b11111111;
		16'b0011000101100001: data <= 8'b11111111;
		16'b0011000111111110: data <= 8'b11111111;
		16'b0011000111111111: data <= 8'b11111111;
		16'b0011001000000000: data <= 8'b11111111;
		16'b0011001000000001: data <= 8'b11111111;
		16'b0011001001001110: data <= 8'b11111111;
		16'b0011001001001111: data <= 8'b11111111;
		16'b0011001001010000: data <= 8'b11111111;
		16'b0011001001010001: data <= 8'b11111111;
		16'b0011001011101110: data <= 8'b11111111;
		16'b0011001011101111: data <= 8'b11111111;
		16'b0011001011110000: data <= 8'b11111111;
		16'b0011001011110001: data <= 8'b11111111;
		16'b0011001100111110: data <= 8'b11111111;
		16'b0011001100111111: data <= 8'b11111111;
		16'b0011001101000000: data <= 8'b11111111;
		16'b0011001101000001: data <= 8'b11111111;
		16'b0011001111011110: data <= 8'b11111111;
		16'b0011001111011111: data <= 8'b11111111;
		16'b0011001111100000: data <= 8'b11111111;
		16'b0011001111100001: data <= 8'b11111111;
		16'b0011010000101110: data <= 8'b11111111;
		16'b0011010000101111: data <= 8'b11111111;
		16'b0011010000110000: data <= 8'b11111111;
		16'b0011010000110001: data <= 8'b11111111;
		16'b0011010011001110: data <= 8'b11111111;
		16'b0011010011001111: data <= 8'b11111111;
		16'b0011010011010000: data <= 8'b11111111;
		16'b0011010011010001: data <= 8'b11111111;
		16'b0011010100011110: data <= 8'b11111111;
		16'b0011010100011111: data <= 8'b11111111;
		16'b0011010100100000: data <= 8'b11111111;
		16'b0011010100100001: data <= 8'b11111111;
		16'b0011010110111110: data <= 8'b11111111;
		16'b0011010110111111: data <= 8'b11111111;
		16'b0011010111000000: data <= 8'b11111111;
		16'b0011010111000001: data <= 8'b11111111;
		16'b0011011000001110: data <= 8'b11111111;
		16'b0011011000001111: data <= 8'b11111111;
		16'b0011011000010000: data <= 8'b11111111;
		16'b0011011000010001: data <= 8'b11111111;
		16'b0011011010101110: data <= 8'b11111111;
		16'b0011011010101111: data <= 8'b11111111;
		16'b0011011010110000: data <= 8'b11111111;
		16'b0011011010110001: data <= 8'b11111111;
		16'b0011011011111110: data <= 8'b11111111;
		16'b0011011011111111: data <= 8'b11111111;
		16'b0011011100000000: data <= 8'b11111111;
		16'b0011011100000001: data <= 8'b11111111;
		16'b0011011110011110: data <= 8'b11111111;
		16'b0011011110011111: data <= 8'b11111111;
		16'b0011011110100000: data <= 8'b11111111;
		16'b0011011110100001: data <= 8'b11111111;
		16'b0011011111101110: data <= 8'b11111111;
		16'b0011011111101111: data <= 8'b11111111;
		16'b0011011111110000: data <= 8'b11111111;
		16'b0011011111110001: data <= 8'b11111111;
		16'b0011100010001110: data <= 8'b11111111;
		16'b0011100010001111: data <= 8'b11111111;
		16'b0011100010010000: data <= 8'b11111111;
		16'b0011100010010001: data <= 8'b11111111;
		16'b0011100011011110: data <= 8'b11111111;
		16'b0011100011011111: data <= 8'b11111111;
		16'b0011100011100000: data <= 8'b11111111;
		16'b0011100011100001: data <= 8'b11111111;
		16'b0011100101111110: data <= 8'b11111111;
		16'b0011100101111111: data <= 8'b11111111;
		16'b0011100110000000: data <= 8'b11111111;
		16'b0011100110000001: data <= 8'b11111111;
		16'b0011100111001110: data <= 8'b11111111;
		16'b0011100111001111: data <= 8'b11111111;
		16'b0011100111010000: data <= 8'b11111111;
		16'b0011100111010001: data <= 8'b11111111;
		16'b0011101001101110: data <= 8'b11111111;
		16'b0011101001101111: data <= 8'b11111111;
		16'b0011101001110000: data <= 8'b11111111;
		16'b0011101001110001: data <= 8'b11111111;
		16'b0011101010111110: data <= 8'b11111111;
		16'b0011101010111111: data <= 8'b11111111;
		16'b0011101011000000: data <= 8'b11111111;
		16'b0011101011000001: data <= 8'b11111111;
		16'b0011101101011110: data <= 8'b11111111;
		16'b0011101101011111: data <= 8'b11111111;
		16'b0011101101100000: data <= 8'b11111111;
		16'b0011101101100001: data <= 8'b11111111;
		16'b0011101110101110: data <= 8'b11111111;
		16'b0011101110101111: data <= 8'b11111111;
		16'b0011101110110000: data <= 8'b11111111;
		16'b0011101110110001: data <= 8'b11111111;
		16'b0011110001001110: data <= 8'b11111111;
		16'b0011110001001111: data <= 8'b11111111;
		16'b0011110001010000: data <= 8'b11111111;
		16'b0011110001010001: data <= 8'b11111111;
		16'b0011110010011110: data <= 8'b11111111;
		16'b0011110010011111: data <= 8'b11111111;
		16'b0011110010100000: data <= 8'b11111111;
		16'b0011110010100001: data <= 8'b11111111;
		16'b0011110100111110: data <= 8'b11111111;
		16'b0011110100111111: data <= 8'b11111111;
		16'b0011110101000000: data <= 8'b11111111;
		16'b0011110101000001: data <= 8'b11111111;
		16'b0011110110001110: data <= 8'b11111111;
		16'b0011110110001111: data <= 8'b11111111;
		16'b0011110110010000: data <= 8'b11111111;
		16'b0011110110010001: data <= 8'b11111111;
		16'b0011111000101110: data <= 8'b11111111;
		16'b0011111000101111: data <= 8'b11111111;
		16'b0011111000110000: data <= 8'b11111111;
		16'b0011111000110001: data <= 8'b11111111;
		16'b0011111001111110: data <= 8'b11111111;
		16'b0011111001111111: data <= 8'b11111111;
		16'b0011111010000000: data <= 8'b11111111;
		16'b0011111010000001: data <= 8'b11111111;
		16'b0011111100011110: data <= 8'b11111111;
		16'b0011111100011111: data <= 8'b11111111;
		16'b0011111100100000: data <= 8'b11111111;
		16'b0011111100100001: data <= 8'b11111111;
		16'b0011111101101110: data <= 8'b11111111;
		16'b0011111101101111: data <= 8'b11111111;
		16'b0011111101110000: data <= 8'b11111111;
		16'b0011111101110001: data <= 8'b11111111;
		16'b0100000000001110: data <= 8'b11111111;
		16'b0100000000001111: data <= 8'b11111111;
		16'b0100000000010000: data <= 8'b11111111;
		16'b0100000000010001: data <= 8'b11111111;
		16'b0100000001011110: data <= 8'b11111111;
		16'b0100000001011111: data <= 8'b11111111;
		16'b0100000001100000: data <= 8'b11111111;
		16'b0100000001100001: data <= 8'b11111111;
		16'b0100000011111110: data <= 8'b11111111;
		16'b0100000011111111: data <= 8'b11111111;
		16'b0100000100000000: data <= 8'b11111111;
		16'b0100000100000001: data <= 8'b11111111;
		16'b0100000101001110: data <= 8'b11111111;
		16'b0100000101001111: data <= 8'b11111111;
		16'b0100000101010000: data <= 8'b11111111;
		16'b0100000101010001: data <= 8'b11111111;
		16'b0100000111101110: data <= 8'b11111111;
		16'b0100000111101111: data <= 8'b11111111;
		16'b0100000111110000: data <= 8'b11111111;
		16'b0100000111110001: data <= 8'b11111111;
		16'b0100001000111110: data <= 8'b11111111;
		16'b0100001000111111: data <= 8'b11111111;
		16'b0100001001000000: data <= 8'b11111111;
		16'b0100001001000001: data <= 8'b11111111;
		16'b0100001011011110: data <= 8'b11111111;
		16'b0100001011011111: data <= 8'b11111111;
		16'b0100001011100000: data <= 8'b11111111;
		16'b0100001011100001: data <= 8'b11111111;
		16'b0100001100101110: data <= 8'b11111111;
		16'b0100001100101111: data <= 8'b11111111;
		16'b0100001100110000: data <= 8'b11111111;
		16'b0100001100110001: data <= 8'b11111111;
		16'b0100001111001110: data <= 8'b11111111;
		16'b0100001111001111: data <= 8'b11111111;
		16'b0100001111010000: data <= 8'b11111111;
		16'b0100001111010001: data <= 8'b11111111;
		16'b0100010000011110: data <= 8'b11111111;
		16'b0100010000011111: data <= 8'b11111111;
		16'b0100010000100000: data <= 8'b11111111;
		16'b0100010000100001: data <= 8'b11111111;
		16'b0100010010111110: data <= 8'b11111111;
		16'b0100010010111111: data <= 8'b11111111;
		16'b0100010011000000: data <= 8'b11111111;
		16'b0100010011000001: data <= 8'b11111111;
		16'b0100010100001110: data <= 8'b11111111;
		16'b0100010100001111: data <= 8'b11111111;
		16'b0100010100010000: data <= 8'b11111111;
		16'b0100010100010001: data <= 8'b11111111;
		16'b0100010110101110: data <= 8'b11111111;
		16'b0100010110101111: data <= 8'b11111111;
		16'b0100010110110000: data <= 8'b11111111;
		16'b0100010110110001: data <= 8'b11111111;
		16'b0100010111111110: data <= 8'b11111111;
		16'b0100010111111111: data <= 8'b11111111;
		16'b0100011000000000: data <= 8'b11111111;
		16'b0100011000000001: data <= 8'b11111111;
		16'b0100011010011110: data <= 8'b11111111;
		16'b0100011010011111: data <= 8'b11111111;
		16'b0100011010100000: data <= 8'b11111111;
		16'b0100011010100001: data <= 8'b11111111;
		16'b0100011011101110: data <= 8'b11111111;
		16'b0100011011101111: data <= 8'b11111111;
		16'b0100011011110000: data <= 8'b11111111;
		16'b0100011011110001: data <= 8'b11111111;
		16'b0100011110001110: data <= 8'b11111111;
		16'b0100011110001111: data <= 8'b11111111;
		16'b0100011110010000: data <= 8'b11111111;
		16'b0100011110010001: data <= 8'b11111111;
		16'b0100011111011110: data <= 8'b11111111;
		16'b0100011111011111: data <= 8'b11111111;
		16'b0100011111100000: data <= 8'b11111111;
		16'b0100011111100001: data <= 8'b11111111;
		16'b0100100001111110: data <= 8'b11111111;
		16'b0100100001111111: data <= 8'b11111111;
		16'b0100100010000000: data <= 8'b11111111;
		16'b0100100010000001: data <= 8'b11111111;
		16'b0100100011001110: data <= 8'b11111111;
		16'b0100100011001111: data <= 8'b11111111;
		16'b0100100011010000: data <= 8'b11111111;
		16'b0100100011010001: data <= 8'b11111111;
		16'b0100100100100000: data <= 8'b11111111;
		16'b0100100100100001: data <= 8'b11111111;
		16'b0100100100100010: data <= 8'b11111111;
		16'b0100100100100011: data <= 8'b11111111;
		16'b0100100100100100: data <= 8'b11111111;
		16'b0100100100100101: data <= 8'b11111111;
		16'b0100100100100110: data <= 8'b11111111;
		16'b0100100100100111: data <= 8'b11111111;
		16'b0100100100101000: data <= 8'b11111111;
		16'b0100100100101001: data <= 8'b11111111;
		16'b0100100100101010: data <= 8'b11111111;
		16'b0100100100101011: data <= 8'b11111111;
		16'b0100100100101100: data <= 8'b11111111;
		16'b0100100100101101: data <= 8'b11111111;
		16'b0100100100101110: data <= 8'b11111111;
		16'b0100100100101111: data <= 8'b11111111;
		16'b0100100100110000: data <= 8'b11111111;
		16'b0100100100110001: data <= 8'b11111111;
		16'b0100100100110010: data <= 8'b11111111;
		16'b0100100100110011: data <= 8'b11111111;
		16'b0100100100110100: data <= 8'b11111111;
		16'b0100100100110101: data <= 8'b11111111;
		16'b0100100100110110: data <= 8'b11111111;
		16'b0100100100110111: data <= 8'b11111111;
		16'b0100100100111000: data <= 8'b11111111;
		16'b0100100100111001: data <= 8'b11111111;
		16'b0100100100111010: data <= 8'b11111111;
		16'b0100100100111011: data <= 8'b11111111;
		16'b0100100100111100: data <= 8'b11111111;
		16'b0100100100111101: data <= 8'b11111111;
		16'b0100100100111110: data <= 8'b11111111;
		16'b0100100100111111: data <= 8'b11111111;
		16'b0100100101000000: data <= 8'b11111111;
		16'b0100100101000001: data <= 8'b11111111;
		16'b0100100101000010: data <= 8'b11111111;
		16'b0100100101000011: data <= 8'b11111111;
		16'b0100100101000100: data <= 8'b11111111;
		16'b0100100101000101: data <= 8'b11111111;
		16'b0100100101000110: data <= 8'b11111111;
		16'b0100100101000111: data <= 8'b11111111;
		16'b0100100101001000: data <= 8'b11111111;
		16'b0100100101001001: data <= 8'b11111111;
		16'b0100100101001010: data <= 8'b11111111;
		16'b0100100101001011: data <= 8'b11111111;
		16'b0100100101001100: data <= 8'b11111111;
		16'b0100100101001101: data <= 8'b11111111;
		16'b0100100101001110: data <= 8'b11111111;
		16'b0100100101001111: data <= 8'b11111111;
		16'b0100100101010000: data <= 8'b11111111;
		16'b0100100101010001: data <= 8'b11111111;
		16'b0100100101010010: data <= 8'b11111111;
		16'b0100100101010011: data <= 8'b11111111;
		16'b0100100101010100: data <= 8'b11111111;
		16'b0100100101010101: data <= 8'b11111111;
		16'b0100100101010110: data <= 8'b11111111;
		16'b0100100101010111: data <= 8'b11111111;
		16'b0100100101011000: data <= 8'b11111111;
		16'b0100100101011001: data <= 8'b11111111;
		16'b0100100101011010: data <= 8'b11111111;
		16'b0100100101011011: data <= 8'b11111111;
		16'b0100100101011100: data <= 8'b11111111;
		16'b0100100101011101: data <= 8'b11111111;
		16'b0100100101011110: data <= 8'b11111111;
		16'b0100100101011111: data <= 8'b11111111;
		16'b0100100101100000: data <= 8'b11111111;
		16'b0100100101100001: data <= 8'b11111111;
		16'b0100100101100010: data <= 8'b11111111;
		16'b0100100101100011: data <= 8'b11111111;
		16'b0100100101100100: data <= 8'b11111111;
		16'b0100100101100101: data <= 8'b11111111;
		16'b0100100101100110: data <= 8'b11111111;
		16'b0100100101100111: data <= 8'b11111111;
		16'b0100100101101000: data <= 8'b11111111;
		16'b0100100101101001: data <= 8'b11111111;
		16'b0100100101101010: data <= 8'b11111111;
		16'b0100100101101011: data <= 8'b11111111;
		16'b0100100101101100: data <= 8'b11111111;
		16'b0100100101101101: data <= 8'b11111111;
		16'b0100100101101110: data <= 8'b11111111;
		16'b0100100101101111: data <= 8'b11111111;
		16'b0100100101110000: data <= 8'b11111111;
		16'b0100100101110001: data <= 8'b11111111;
		16'b0100100101110010: data <= 8'b11111111;
		16'b0100100101110011: data <= 8'b11111111;
		16'b0100100101110100: data <= 8'b11111111;
		16'b0100100101110101: data <= 8'b11111111;
		16'b0100100101110110: data <= 8'b11111111;
		16'b0100100101110111: data <= 8'b11111111;
		16'b0100100101111000: data <= 8'b11111111;
		16'b0100100101111001: data <= 8'b11111111;
		16'b0100100101111010: data <= 8'b11111111;
		16'b0100100101111011: data <= 8'b11111111;
		16'b0100100101111100: data <= 8'b11111111;
		16'b0100100101111101: data <= 8'b11111111;
		16'b0100100101111110: data <= 8'b11111111;
		16'b0100100101111111: data <= 8'b11111111;
		16'b0100100110000000: data <= 8'b11111111;
		16'b0100100110000001: data <= 8'b11111111;
		16'b0100100110000010: data <= 8'b11111111;
		16'b0100100110000011: data <= 8'b11111111;
		16'b0100100110000100: data <= 8'b11111111;
		16'b0100100110000101: data <= 8'b11111111;
		16'b0100100110000110: data <= 8'b11111111;
		16'b0100100110000111: data <= 8'b11111111;
		16'b0100100110001000: data <= 8'b11111111;
		16'b0100100110001001: data <= 8'b11111111;
		16'b0100100110001010: data <= 8'b11111111;
		16'b0100100110001011: data <= 8'b11111111;
		16'b0100100110001100: data <= 8'b11111111;
		16'b0100100110001101: data <= 8'b11111111;
		16'b0100100110001110: data <= 8'b11111111;
		16'b0100100110001111: data <= 8'b11111111;
		16'b0100100110010000: data <= 8'b11111111;
		16'b0100100110010001: data <= 8'b11111111;
		16'b0100100110010010: data <= 8'b11111111;
		16'b0100100110010011: data <= 8'b11111111;
		16'b0100100110010100: data <= 8'b11111111;
		16'b0100100110010101: data <= 8'b11111111;
		16'b0100100110010110: data <= 8'b11111111;
		16'b0100100110010111: data <= 8'b11111111;
		16'b0100100110011000: data <= 8'b11111111;
		16'b0100100110011001: data <= 8'b11111111;
		16'b0100100110011010: data <= 8'b11111111;
		16'b0100100110011011: data <= 8'b11111111;
		16'b0100100110011100: data <= 8'b11111111;
		16'b0100100110011101: data <= 8'b11111111;
		16'b0100100110011110: data <= 8'b11111111;
		16'b0100100110011111: data <= 8'b11111111;
		16'b0100100110100000: data <= 8'b11111111;
		16'b0100100110100001: data <= 8'b11111111;
		16'b0100100110100010: data <= 8'b11111111;
		16'b0100100110100011: data <= 8'b11111111;
		16'b0100100110100100: data <= 8'b11111111;
		16'b0100100110100101: data <= 8'b11111111;
		16'b0100100110100110: data <= 8'b11111111;
		16'b0100100110100111: data <= 8'b11111111;
		16'b0100100110101000: data <= 8'b11111111;
		16'b0100100110101001: data <= 8'b11111111;
		16'b0100100110101010: data <= 8'b11111111;
		16'b0100100110101011: data <= 8'b11111111;
		16'b0100100110101100: data <= 8'b11111111;
		16'b0100100110101101: data <= 8'b11111111;
		16'b0100100110101110: data <= 8'b11111111;
		16'b0100100110101111: data <= 8'b11111111;
		16'b0100100110110000: data <= 8'b11111111;
		16'b0100100110110001: data <= 8'b11111111;
		16'b0100100110110010: data <= 8'b11111111;
		16'b0100100110110011: data <= 8'b11111111;
		16'b0100100110110100: data <= 8'b11111111;
		16'b0100100110110101: data <= 8'b11111111;
		16'b0100100110110110: data <= 8'b11111111;
		16'b0100100110110111: data <= 8'b11111111;
		16'b0100100110111000: data <= 8'b11111111;
		16'b0100100110111001: data <= 8'b11111111;
		16'b0100100110111010: data <= 8'b11111111;
		16'b0100100110111011: data <= 8'b11111111;
		16'b0100100110111100: data <= 8'b11111111;
		16'b0100100110111101: data <= 8'b11111111;
		16'b0100100110111110: data <= 8'b11111111;
		16'b0100100110111111: data <= 8'b11111111;
		16'b0100100111000000: data <= 8'b11111111;
		16'b0100100111000001: data <= 8'b11111111;
		16'b0100100111000010: data <= 8'b11111111;
		16'b0100100111000011: data <= 8'b11111111;
		16'b0100100111000100: data <= 8'b11111111;
		16'b0100100111000101: data <= 8'b11111111;
		16'b0100100111000110: data <= 8'b11111111;
		16'b0100100111000111: data <= 8'b11111111;
		16'b0100100111001000: data <= 8'b11111111;
		16'b0100100111001001: data <= 8'b11111111;
		16'b0100100111001010: data <= 8'b11111111;
		16'b0100100111001011: data <= 8'b11111111;
		16'b0100100111001100: data <= 8'b11111111;
		16'b0100100111001101: data <= 8'b11111111;
		16'b0100100111001110: data <= 8'b11111111;
		16'b0100100111001111: data <= 8'b11111111;
		16'b0100100111010000: data <= 8'b11111111;
		16'b0100100111010001: data <= 8'b11111111;
		16'b0100100111010010: data <= 8'b11111111;
		16'b0100100111010011: data <= 8'b11111111;
		16'b0100100111010100: data <= 8'b11111111;
		16'b0100100111010101: data <= 8'b11111111;
		16'b0100100111010110: data <= 8'b11111111;
		16'b0100100111010111: data <= 8'b11111111;
		16'b0100100111011000: data <= 8'b11111111;
		16'b0100100111011001: data <= 8'b11111111;
		16'b0100100111011010: data <= 8'b11111111;
		16'b0100100111011011: data <= 8'b11111111;
		16'b0100100111011100: data <= 8'b11111111;
		16'b0100100111011101: data <= 8'b11111111;
		16'b0100100111011110: data <= 8'b11111111;
		16'b0100100111011111: data <= 8'b11111111;
		16'b0100100111100000: data <= 8'b11111111;
		16'b0100100111100001: data <= 8'b11111111;
		16'b0100100111100010: data <= 8'b11111111;
		16'b0100100111100011: data <= 8'b11111111;
		16'b0100100111100100: data <= 8'b11111111;
		16'b0100100111100101: data <= 8'b11111111;
		16'b0100100111100110: data <= 8'b11111111;
		16'b0100100111100111: data <= 8'b11111111;
		16'b0100100111101000: data <= 8'b11111111;
		16'b0100100111101001: data <= 8'b11111111;
		16'b0100100111101010: data <= 8'b11111111;
		16'b0100100111101011: data <= 8'b11111111;
		16'b0100100111101100: data <= 8'b11111111;
		16'b0100100111101101: data <= 8'b11111111;
		16'b0100100111101110: data <= 8'b11111111;
		16'b0100100111101111: data <= 8'b11111111;
		16'b0100100111110000: data <= 8'b11111111;
		16'b0100100111110001: data <= 8'b11111111;
		16'b0100100111110010: data <= 8'b11111111;
		16'b0100100111110011: data <= 8'b11111111;
		16'b0100100111110100: data <= 8'b11111111;
		16'b0100100111110101: data <= 8'b11111111;
		16'b0100100111110110: data <= 8'b11111111;
		16'b0100100111110111: data <= 8'b11111111;
		16'b0100100111111000: data <= 8'b11111111;
		16'b0100100111111001: data <= 8'b11111111;
		16'b0100100111111010: data <= 8'b11111111;
		16'b0100100111111011: data <= 8'b11111111;
		16'b0100100111111100: data <= 8'b11111111;
		16'b0100100111111101: data <= 8'b11111111;
		16'b0100100111111110: data <= 8'b11111111;
		16'b0100100111111111: data <= 8'b11111111;
		16'b0100101000000000: data <= 8'b11111111;
		16'b0100101000000001: data <= 8'b11111111;
		16'b0100101000000010: data <= 8'b11111111;
		16'b0100101000000011: data <= 8'b11111111;
		16'b0100101000000100: data <= 8'b11111111;
		16'b0100101000000101: data <= 8'b11111111;
		16'b0100101000000110: data <= 8'b11111111;
		16'b0100101000000111: data <= 8'b11111111;
		16'b0100101000001000: data <= 8'b11111111;
		16'b0100101000001001: data <= 8'b11111111;
		16'b0100101000001010: data <= 8'b11111111;
		16'b0100101000001011: data <= 8'b11111111;
		16'b0100101000001100: data <= 8'b11111111;
		16'b0100101000001101: data <= 8'b11111111;
		16'b0100101000001110: data <= 8'b11111111;
		16'b0100101000001111: data <= 8'b11111111;
		16'b0100101000010000: data <= 8'b11111111;
		16'b0100101000010001: data <= 8'b11111111;
		16'b0100101000010010: data <= 8'b11111111;
		16'b0100101000010011: data <= 8'b11111111;
		16'b0100101000010100: data <= 8'b11111111;
		16'b0100101000010101: data <= 8'b11111111;
		16'b0100101000010110: data <= 8'b11111111;
		16'b0100101000010111: data <= 8'b11111111;
		16'b0100101000011000: data <= 8'b11111111;
		16'b0100101000011001: data <= 8'b11111111;
		16'b0100101000011010: data <= 8'b11111111;
		16'b0100101000011011: data <= 8'b11111111;
		16'b0100101000011100: data <= 8'b11111111;
		16'b0100101000011101: data <= 8'b11111111;
		16'b0100101000011110: data <= 8'b11111111;
		16'b0100101000011111: data <= 8'b11111111;
		16'b0100101000100000: data <= 8'b11111111;
		16'b0100101000100001: data <= 8'b11111111;
		16'b0100101000100010: data <= 8'b11111111;
		16'b0100101000100011: data <= 8'b11111111;
		16'b0100101000100100: data <= 8'b11111111;
		16'b0100101000100101: data <= 8'b11111111;
		16'b0100101000100110: data <= 8'b11111111;
		16'b0100101000100111: data <= 8'b11111111;
		16'b0100101000101000: data <= 8'b11111111;
		16'b0100101000101001: data <= 8'b11111111;
		16'b0100101000101010: data <= 8'b11111111;
		16'b0100101000101011: data <= 8'b11111111;
		16'b0100101000101100: data <= 8'b11111111;
		16'b0100101000101101: data <= 8'b11111111;
		16'b0100101000101110: data <= 8'b11111111;
		16'b0100101000101111: data <= 8'b11111111;
		16'b0100101000110000: data <= 8'b11111111;
		16'b0100101000110001: data <= 8'b11111111;
		16'b0100101000110010: data <= 8'b11111111;
		16'b0100101000110011: data <= 8'b11111111;
		16'b0100101000110100: data <= 8'b11111111;
		16'b0100101000110101: data <= 8'b11111111;
		16'b0100101000110110: data <= 8'b11111111;
		16'b0100101000110111: data <= 8'b11111111;
		16'b0100101000111000: data <= 8'b11111111;
		16'b0100101000111001: data <= 8'b11111111;
		16'b0100101000111010: data <= 8'b11111111;
		16'b0100101000111011: data <= 8'b11111111;
		16'b0100101000111100: data <= 8'b11111111;
		16'b0100101000111101: data <= 8'b11111111;
		16'b0100101000111110: data <= 8'b11111111;
		16'b0100101000111111: data <= 8'b11111111;
		16'b0100101001000000: data <= 8'b11111111;
		16'b0100101001000001: data <= 8'b11111111;
		16'b0100101001000010: data <= 8'b11111111;
		16'b0100101001000011: data <= 8'b11111111;
		16'b0100101001000100: data <= 8'b11111111;
		16'b0100101001000101: data <= 8'b11111111;
		16'b0100101001000110: data <= 8'b11111111;
		16'b0100101001000111: data <= 8'b11111111;
		16'b0100101001001000: data <= 8'b11111111;
		16'b0100101001001001: data <= 8'b11111111;
		16'b0100101001001010: data <= 8'b11111111;
		16'b0100101001001011: data <= 8'b11111111;
		16'b0100101001001100: data <= 8'b11111111;
		16'b0100101001001101: data <= 8'b11111111;
		16'b0100101001001110: data <= 8'b11111111;
		16'b0100101001001111: data <= 8'b11111111;
		16'b0100101001010000: data <= 8'b11111111;
		16'b0100101001010001: data <= 8'b11111111;
		16'b0100101001010010: data <= 8'b11111111;
		16'b0100101001010011: data <= 8'b11111111;
		16'b0100101001010100: data <= 8'b11111111;
		16'b0100101001010101: data <= 8'b11111111;
		16'b0100101001010110: data <= 8'b11111111;
		16'b0100101001010111: data <= 8'b11111111;
		16'b0100101001011000: data <= 8'b11111111;
		16'b0100101001011001: data <= 8'b11111111;
		16'b0100101001011010: data <= 8'b11111111;
		16'b0100101001011011: data <= 8'b11111111;
		16'b0100101001011100: data <= 8'b11111111;
		16'b0100101001011101: data <= 8'b11111111;
		16'b0100101001011110: data <= 8'b11111111;
		16'b0100101001011111: data <= 8'b11111111;
		16'b0100101001100000: data <= 8'b11111111;
		16'b0100101001100001: data <= 8'b11111111;
		16'b0100101001100010: data <= 8'b11111111;
		16'b0100101001100011: data <= 8'b11111111;
		16'b0100101001100100: data <= 8'b11111111;
		16'b0100101001100101: data <= 8'b11111111;
		16'b0100101001100110: data <= 8'b11111111;
		16'b0100101001100111: data <= 8'b11111111;
		16'b0100101001101000: data <= 8'b11111111;
		16'b0100101001101001: data <= 8'b11111111;
		16'b0100101001101010: data <= 8'b11111111;
		16'b0100101001101011: data <= 8'b11111111;
		16'b0100101001101100: data <= 8'b11111111;
		16'b0100101001101101: data <= 8'b11111111;
		16'b0100101001101110: data <= 8'b11111111;
		16'b0100101001101111: data <= 8'b11111111;
		16'b0100101001110000: data <= 8'b11111111;
		16'b0100101001110001: data <= 8'b11111111;
		16'b0100101001110010: data <= 8'b11111111;
		16'b0100101001110011: data <= 8'b11111111;
		16'b0100101001110100: data <= 8'b11111111;
		16'b0100101001110101: data <= 8'b11111111;
		16'b0100101001110110: data <= 8'b11111111;
		16'b0100101001110111: data <= 8'b11111111;
		16'b0100101001111000: data <= 8'b11111111;
		16'b0100101001111001: data <= 8'b11111111;
		16'b0100101001111010: data <= 8'b11111111;
		16'b0100101001111011: data <= 8'b11111111;
		16'b0100101001111100: data <= 8'b11111111;
		16'b0100101001111101: data <= 8'b11111111;
		16'b0100101001111110: data <= 8'b11111111;
		16'b0100101001111111: data <= 8'b11111111;
		16'b0100101010000000: data <= 8'b11111111;
		16'b0100101010000001: data <= 8'b11111111;
		16'b0100101010000010: data <= 8'b11111111;
		16'b0100101010000011: data <= 8'b11111111;
		16'b0100101010000100: data <= 8'b11111111;
		16'b0100101010000101: data <= 8'b11111111;
		16'b0100101010000110: data <= 8'b11111111;
		16'b0100101010000111: data <= 8'b11111111;
		16'b0100101010001000: data <= 8'b11111111;
		16'b0100101010001001: data <= 8'b11111111;
		16'b0100101010001010: data <= 8'b11111111;
		16'b0100101010001011: data <= 8'b11111111;
		16'b0100101010001100: data <= 8'b11111111;
		16'b0100101010001101: data <= 8'b11111111;
		16'b0100101010001110: data <= 8'b11111111;
		16'b0100101010001111: data <= 8'b11111111;
		16'b0100101010010000: data <= 8'b11111111;
		16'b0100101010010001: data <= 8'b11111111;
		16'b0100101010010010: data <= 8'b11111111;
		16'b0100101010010011: data <= 8'b11111111;
		16'b0100101010010100: data <= 8'b11111111;
		16'b0100101010010101: data <= 8'b11111111;
		16'b0100101010010110: data <= 8'b11111111;
		16'b0100101010010111: data <= 8'b11111111;
		16'b0100101010011000: data <= 8'b11111111;
		16'b0100101010011001: data <= 8'b11111111;
		16'b0100101010011010: data <= 8'b11111111;
		16'b0100101010011011: data <= 8'b11111111;
		16'b0100101010011100: data <= 8'b11111111;
		16'b0100101010011101: data <= 8'b11111111;
		16'b0100101010011110: data <= 8'b11111111;
		16'b0100101010011111: data <= 8'b11111111;
		16'b0100101010100000: data <= 8'b11111111;
		16'b0100101010100001: data <= 8'b11111111;
		16'b0100101010100010: data <= 8'b11111111;
		16'b0100101010100011: data <= 8'b11111111;
		16'b0100101010100100: data <= 8'b11111111;
		16'b0100101010100101: data <= 8'b11111111;
		16'b0100101010100110: data <= 8'b11111111;
		16'b0100101010100111: data <= 8'b11111111;
		16'b0100101010101000: data <= 8'b11111111;
		16'b0100101010101001: data <= 8'b11111111;
		16'b0100101010101010: data <= 8'b11111111;
		16'b0100101010101011: data <= 8'b11111111;
		16'b0100101010101100: data <= 8'b11111111;
		16'b0100101010101101: data <= 8'b11111111;
		16'b0100101010101110: data <= 8'b11111111;
		16'b0100101010101111: data <= 8'b11111111;
		16'b0100101010110000: data <= 8'b11111111;
		16'b0100101010110001: data <= 8'b11111111;
		16'b0100101010110010: data <= 8'b11111111;
		16'b0100101010110011: data <= 8'b11111111;
		16'b0100101010110100: data <= 8'b11111111;
		16'b0100101010110101: data <= 8'b11111111;
		16'b0100101010110110: data <= 8'b11111111;
		16'b0100101010110111: data <= 8'b11111111;
		16'b0100101010111000: data <= 8'b11111111;
		16'b0100101010111001: data <= 8'b11111111;
		16'b0100101010111010: data <= 8'b11111111;
		16'b0100101010111011: data <= 8'b11111111;
		16'b0100101010111100: data <= 8'b11111111;
		16'b0100101010111101: data <= 8'b11111111;
		16'b0100101010111110: data <= 8'b11111111;
		16'b0100101010111111: data <= 8'b11111111;
		16'b0100101011000000: data <= 8'b11111111;
		16'b0100101011000001: data <= 8'b11111111;
		16'b0100101011000010: data <= 8'b11111111;
		16'b0100101011000011: data <= 8'b11111111;
		16'b0100101011000100: data <= 8'b11111111;
		16'b0100101011000101: data <= 8'b11111111;
		16'b0100101011000110: data <= 8'b11111111;
		16'b0100101011000111: data <= 8'b11111111;
		16'b0100101011001000: data <= 8'b11111111;
		16'b0100101011001001: data <= 8'b11111111;
		16'b0100101011001010: data <= 8'b11111111;
		16'b0100101011001011: data <= 8'b11111111;
		16'b0100101011001100: data <= 8'b11111111;
		16'b0100101011001101: data <= 8'b11111111;
		16'b0100101011001110: data <= 8'b11111111;
		16'b0100101011001111: data <= 8'b11111111;
		16'b0100101011010000: data <= 8'b11111111;
		16'b0100101011010001: data <= 8'b11111111;
		16'b0100101011010010: data <= 8'b11111111;
		16'b0100101011010011: data <= 8'b11111111;
		16'b0100101011010100: data <= 8'b11111111;
		16'b0100101011010101: data <= 8'b11111111;
		16'b0100101011010110: data <= 8'b11111111;
		16'b0100101011010111: data <= 8'b11111111;
		16'b0100101011011000: data <= 8'b11111111;
		16'b0100101011011001: data <= 8'b11111111;
		16'b0100101011011010: data <= 8'b11111111;
		16'b0100101011011011: data <= 8'b11111111;
		16'b0100101011011100: data <= 8'b11111111;
		16'b0100101011011101: data <= 8'b11111111;
		16'b0100101011011110: data <= 8'b11111111;
		16'b0100101011011111: data <= 8'b11111111;
		16'b0100101011100000: data <= 8'b11111111;
		16'b0100101011100001: data <= 8'b11111111;
		16'b0100101011100010: data <= 8'b11111111;
		16'b0100101011100011: data <= 8'b11111111;
		16'b0100101011100100: data <= 8'b11111111;
		16'b0100101011100101: data <= 8'b11111111;
		16'b0100101011100110: data <= 8'b11111111;
		16'b0100101011100111: data <= 8'b11111111;
		16'b0100101011101000: data <= 8'b11111111;
		16'b0100101011101001: data <= 8'b11111111;
		16'b0100101011101010: data <= 8'b11111111;
		16'b0100101011101011: data <= 8'b11111111;
		16'b0100101011101100: data <= 8'b11111111;
		16'b0100101011101101: data <= 8'b11111111;
		16'b0100101011101110: data <= 8'b11111111;
		16'b0100101011101111: data <= 8'b11111111;
		16'b0100101011110000: data <= 8'b11111111;
		16'b0100101011110001: data <= 8'b11111111;
		16'b0100101011110010: data <= 8'b11111111;
		16'b0100101011110011: data <= 8'b11111111;
		16'b0100101011110100: data <= 8'b11111111;
		16'b0100101011110101: data <= 8'b11111111;
		16'b0100101011110110: data <= 8'b11111111;
		16'b0100101011110111: data <= 8'b11111111;
		16'b0100101011111000: data <= 8'b11111111;
		16'b0100101011111001: data <= 8'b11111111;
		16'b0100101011111010: data <= 8'b11111111;
		16'b0100101011111011: data <= 8'b11111111;
		16'b0100101011111100: data <= 8'b11111111;
		16'b0100101011111101: data <= 8'b11111111;
		16'b0100101011111110: data <= 8'b11111111;
		16'b0100101011111111: data <= 8'b11111111;
		16'b0100101100000000: data <= 8'b11111111;
		16'b0100101100000001: data <= 8'b11111111;
		16'b0100101100000010: data <= 8'b11111111;
		16'b0100101100000011: data <= 8'b11111111;
		16'b0100101100000100: data <= 8'b11111111;
		16'b0100101100000101: data <= 8'b11111111;
		16'b0100101100000110: data <= 8'b11111111;
		16'b0100101100000111: data <= 8'b11111111;
		16'b0100101100001000: data <= 8'b11111111;
		16'b0100101100001001: data <= 8'b11111111;
		16'b0100101100001010: data <= 8'b11111111;
		16'b0100101100001011: data <= 8'b11111111;
		16'b0100101100001100: data <= 8'b11111111;
		16'b0100101100001101: data <= 8'b11111111;
		16'b0100101100001110: data <= 8'b11111111;
		16'b0100101100001111: data <= 8'b11111111;
		16'b0100101100010000: data <= 8'b11111111;
		16'b0100101100010001: data <= 8'b11111111;
		16'b0100101100010010: data <= 8'b11111111;
		16'b0100101100010011: data <= 8'b11111111;
		16'b0100101100010100: data <= 8'b11111111;
		16'b0100101100010101: data <= 8'b11111111;
		16'b0100101100010110: data <= 8'b11111111;
		16'b0100101100010111: data <= 8'b11111111;
		16'b0100101100011000: data <= 8'b11111111;
		16'b0100101100011001: data <= 8'b11111111;
		16'b0100101100011010: data <= 8'b11111111;
		16'b0100101100011011: data <= 8'b11111111;
		16'b0100101100011100: data <= 8'b11111111;
		16'b0100101100011101: data <= 8'b11111111;
		16'b0100101100011110: data <= 8'b11111111;
		16'b0100101100011111: data <= 8'b11111111;
		16'b0100101100100000: data <= 8'b11111111;
		16'b0100101100100001: data <= 8'b11111111;
		16'b0100101100100010: data <= 8'b11111111;
		16'b0100101100100011: data <= 8'b11111111;
		16'b0100101100100100: data <= 8'b11111111;
		16'b0100101100100101: data <= 8'b11111111;
		16'b0100101100100110: data <= 8'b11111111;
		16'b0100101100100111: data <= 8'b11111111;
		16'b0100101100101000: data <= 8'b11111111;
		16'b0100101100101001: data <= 8'b11111111;
		16'b0100101100101010: data <= 8'b11111111;
		16'b0100101100101011: data <= 8'b11111111;
		16'b0100101100101100: data <= 8'b11111111;
		16'b0100101100101101: data <= 8'b11111111;
		16'b0100101100101110: data <= 8'b11111111;
		16'b0100101100101111: data <= 8'b11111111;
		16'b0100101100110000: data <= 8'b11111111;
		16'b0100101100110001: data <= 8'b11111111;
		16'b0100101100110010: data <= 8'b11111111;
		16'b0100101100110011: data <= 8'b11111111;
		16'b0100101100110100: data <= 8'b11111111;
		16'b0100101100110101: data <= 8'b11111111;
		16'b0100101100110110: data <= 8'b11111111;
		16'b0100101100110111: data <= 8'b11111111;
		16'b0100101100111000: data <= 8'b11111111;
		16'b0100101100111001: data <= 8'b11111111;
		16'b0100101100111010: data <= 8'b11111111;
		16'b0100101100111011: data <= 8'b11111111;
		16'b0100101100111100: data <= 8'b11111111;
		16'b0100101100111101: data <= 8'b11111111;
		16'b0100101100111110: data <= 8'b11111111;
		16'b0100101100111111: data <= 8'b11111111;
		16'b0100101101000000: data <= 8'b11111111;
		16'b0100101101000001: data <= 8'b11111111;
		16'b0100101101000010: data <= 8'b11111111;
		16'b0100101101000011: data <= 8'b11111111;
		16'b0100101101000100: data <= 8'b11111111;
		16'b0100101101000101: data <= 8'b11111111;
		16'b0100101101000110: data <= 8'b11111111;
		16'b0100101101000111: data <= 8'b11111111;
		16'b0100101101001000: data <= 8'b11111111;
		16'b0100101101001001: data <= 8'b11111111;
		16'b0100101101001010: data <= 8'b11111111;
		16'b0100101101001011: data <= 8'b11111111;
		16'b0100101101001100: data <= 8'b11111111;
		16'b0100101101001101: data <= 8'b11111111;
		16'b0100101101001110: data <= 8'b11111111;
		16'b0100101101001111: data <= 8'b11111111;
		16'b0100101101010000: data <= 8'b11111111;
		16'b0100101101010001: data <= 8'b11111111;
		16'b0100101101010010: data <= 8'b11111111;
		16'b0100101101010011: data <= 8'b11111111;
		16'b0100101101010100: data <= 8'b11111111;
		16'b0100101101010101: data <= 8'b11111111;
		16'b0100101101010110: data <= 8'b11111111;
		16'b0100101101010111: data <= 8'b11111111;
		16'b0100101101011000: data <= 8'b11111111;
		16'b0100101101011001: data <= 8'b11111111;
		16'b0100101101011010: data <= 8'b11111111;
		16'b0100101101011011: data <= 8'b11111111;
		16'b0100101101011100: data <= 8'b11111111;
		16'b0100101101011101: data <= 8'b11111111;
		16'b0100101101011110: data <= 8'b11111111;
		16'b0100101101011111: data <= 8'b11111111;
		16'b0100101101100000: data <= 8'b11111111;
		16'b0100101101100001: data <= 8'b11111111;
		16'b0100101101100010: data <= 8'b11111111;
		16'b0100101101100011: data <= 8'b11111111;
		16'b0100101101100100: data <= 8'b11111111;
		16'b0100101101100101: data <= 8'b11111111;
		16'b0100101101100110: data <= 8'b11111111;
		16'b0100101101100111: data <= 8'b11111111;
		16'b0100101101101000: data <= 8'b11111111;
		16'b0100101101101001: data <= 8'b11111111;
		16'b0100101101101010: data <= 8'b11111111;
		16'b0100101101101011: data <= 8'b11111111;
		16'b0100101101101100: data <= 8'b11111111;
		16'b0100101101101101: data <= 8'b11111111;
		16'b0100101101101110: data <= 8'b11111111;
		16'b0100101101101111: data <= 8'b11111111;
		16'b0100101101110000: data <= 8'b11111111;
		16'b0100101101110001: data <= 8'b11111111;
		16'b0100101101110010: data <= 8'b11111111;
		16'b0100101101110011: data <= 8'b11111111;
		16'b0100101101110100: data <= 8'b11111111;
		16'b0100101101110101: data <= 8'b11111111;
		16'b0100101101110110: data <= 8'b11111111;
		16'b0100101101110111: data <= 8'b11111111;
		16'b0100101101111000: data <= 8'b11111111;
		16'b0100101101111001: data <= 8'b11111111;
		16'b0100101101111010: data <= 8'b11111111;
		16'b0100101101111011: data <= 8'b11111111;
		16'b0100101101111100: data <= 8'b11111111;
		16'b0100101101111101: data <= 8'b11111111;
		16'b0100101101111110: data <= 8'b11111111;
		16'b0100101101111111: data <= 8'b11111111;
		16'b0100101110000000: data <= 8'b11111111;
		16'b0100101110000001: data <= 8'b11111111;
		16'b0100101110000010: data <= 8'b11111111;
		16'b0100101110000011: data <= 8'b11111111;
		16'b0100101110000100: data <= 8'b11111111;
		16'b0100101110000101: data <= 8'b11111111;
		16'b0100101110000110: data <= 8'b11111111;
		16'b0100101110000111: data <= 8'b11111111;
		16'b0100101110001000: data <= 8'b11111111;
		16'b0100101110001001: data <= 8'b11111111;
		16'b0100101110001010: data <= 8'b11111111;
		16'b0100101110001011: data <= 8'b11111111;
		16'b0100101110001100: data <= 8'b11111111;
		16'b0100101110001101: data <= 8'b11111111;
		16'b0100101110001110: data <= 8'b11111111;
		16'b0100101110001111: data <= 8'b11111111;
		16'b0100101110010000: data <= 8'b11111111;
		16'b0100101110010001: data <= 8'b11111111;
		16'b0100101110010010: data <= 8'b11111111;
		16'b0100101110010011: data <= 8'b11111111;
		16'b0100101110010100: data <= 8'b11111111;
		16'b0100101110010101: data <= 8'b11111111;
		16'b0100101110010110: data <= 8'b11111111;
		16'b0100101110010111: data <= 8'b11111111;
		16'b0100101110011000: data <= 8'b11111111;
		16'b0100101110011001: data <= 8'b11111111;
		16'b0100101110011010: data <= 8'b11111111;
		16'b0100101110011011: data <= 8'b11111111;
		16'b0100101110011100: data <= 8'b11111111;
		16'b0100101110011101: data <= 8'b11111111;
		16'b0100101110011110: data <= 8'b11111111;
		16'b0100101110011111: data <= 8'b11111111;
		16'b0100101110100000: data <= 8'b11111111;
		16'b0100101110100001: data <= 8'b11111111;
		16'b0100101110100010: data <= 8'b11111111;
		16'b0100101110100011: data <= 8'b11111111;
		16'b0100101110100100: data <= 8'b11111111;
		16'b0100101110100101: data <= 8'b11111111;
		16'b0100101110100110: data <= 8'b11111111;
		16'b0100101110100111: data <= 8'b11111111;
		16'b0100101110101000: data <= 8'b11111111;
		16'b0100101110101001: data <= 8'b11111111;
		16'b0100101110101010: data <= 8'b11111111;
		16'b0100101110101011: data <= 8'b11111111;
		16'b0100101110101100: data <= 8'b11111111;
		16'b0100101110101101: data <= 8'b11111111;
		16'b0100101110101110: data <= 8'b11111111;
		16'b0100101110101111: data <= 8'b11111111;
		16'b0100101110110000: data <= 8'b11111111;
		16'b0100101110110001: data <= 8'b11111111;
		16'b0100101110110010: data <= 8'b11111111;
		16'b0100101110110011: data <= 8'b11111111;
		16'b0100101110110100: data <= 8'b11111111;
		16'b0100101110110101: data <= 8'b11111111;
		16'b0100101110110110: data <= 8'b11111111;
		16'b0100101110110111: data <= 8'b11111111;
		16'b0100101110111000: data <= 8'b11111111;
		16'b0100101110111001: data <= 8'b11111111;
		16'b0100101110111010: data <= 8'b11111111;
		16'b0100101110111011: data <= 8'b11111111;
		16'b0100101110111100: data <= 8'b11111111;
		16'b0100101110111101: data <= 8'b11111111;
		16'b0100101110111110: data <= 8'b11111111;
		16'b0100101110111111: data <= 8'b11111111;
		16'b0100101111000000: data <= 8'b11111111;
		16'b0100101111000001: data <= 8'b11111111;
		16'b0100101111000010: data <= 8'b11111111;
		16'b0100101111000011: data <= 8'b11111111;
		16'b0100101111000100: data <= 8'b11111111;
		16'b0100101111000101: data <= 8'b11111111;
		16'b0100101111000110: data <= 8'b11111111;
		16'b0100101111000111: data <= 8'b11111111;
		16'b0100101111001000: data <= 8'b11111111;
		16'b0100101111001001: data <= 8'b11111111;
		16'b0100101111001010: data <= 8'b11111111;
		16'b0100101111001011: data <= 8'b11111111;
		16'b0100101111001100: data <= 8'b11111111;
		16'b0100101111001101: data <= 8'b11111111;
		16'b0100101111001110: data <= 8'b11111111;
		16'b0100101111001111: data <= 8'b11111111;
		16'b0100101111010000: data <= 8'b11111111;
		16'b0100101111010001: data <= 8'b11111111;
		16'b0100101111010010: data <= 8'b11111111;
		16'b0100101111010011: data <= 8'b11111111;
		16'b0100101111010100: data <= 8'b11111111;
		16'b0100101111010101: data <= 8'b11111111;
		16'b0100101111010110: data <= 8'b11111111;
		16'b0100101111010111: data <= 8'b11111111;
		16'b0100101111011000: data <= 8'b11111111;
		16'b0100101111011001: data <= 8'b11111111;
		16'b0100101111011010: data <= 8'b11111111;
		16'b0100101111011011: data <= 8'b11111111;
		16'b0100101111011100: data <= 8'b11111111;
		16'b0100101111011101: data <= 8'b11111111;
		16'b0100101111011110: data <= 8'b11111111;
		16'b0100101111011111: data <= 8'b11111111;
		16'b0100101111100000: data <= 8'b11111111;
		16'b0100101111100001: data <= 8'b11111111;
		16'b0100101111100010: data <= 8'b11111111;
		16'b0100101111100011: data <= 8'b11111111;
		16'b0100101111100100: data <= 8'b11111111;
		16'b0100101111100101: data <= 8'b11111111;
		16'b0100101111100110: data <= 8'b11111111;
		16'b0100101111100111: data <= 8'b11111111;
		16'b0100101111101000: data <= 8'b11111111;
		16'b0100101111101001: data <= 8'b11111111;
		16'b0100101111101010: data <= 8'b11111111;
		16'b0100101111101011: data <= 8'b11111111;
		16'b0100101111101100: data <= 8'b11111111;
		16'b0100101111101101: data <= 8'b11111111;
		16'b0100101111101110: data <= 8'b11111111;
		16'b0100101111101111: data <= 8'b11111111;
		16'b0100101111110000: data <= 8'b11111111;
		16'b0100101111110001: data <= 8'b11111111;
		16'b0100101111110010: data <= 8'b11111111;
		16'b0100101111110011: data <= 8'b11111111;
		16'b0100101111110100: data <= 8'b11111111;
		16'b0100101111110101: data <= 8'b11111111;
		16'b0100101111110110: data <= 8'b11111111;
		16'b0100101111110111: data <= 8'b11111111;
		16'b0100101111111000: data <= 8'b11111111;
		16'b0100101111111001: data <= 8'b11111111;
		16'b0100101111111010: data <= 8'b11111111;
		16'b0100101111111011: data <= 8'b11111111;
		16'b0100101111111100: data <= 8'b11111111;
		16'b0100101111111101: data <= 8'b11111111;
		16'b0100101111111110: data <= 8'b11111111;
		16'b0100101111111111: data <= 8'b11111111;
		16'b0100110000000000: data <= 8'b11111111;
		16'b0100110000000001: data <= 8'b11111111;
		16'b0100110000000010: data <= 8'b11111111;
		16'b0100110000000011: data <= 8'b11111111;
		16'b0100110000000100: data <= 8'b11111111;
		16'b0100110000000101: data <= 8'b11111111;
		16'b0100110000000110: data <= 8'b11111111;
		16'b0100110000000111: data <= 8'b11111111;
		16'b0100110000001000: data <= 8'b11111111;
		16'b0100110000001001: data <= 8'b11111111;
		16'b0100110000001010: data <= 8'b11111111;
		16'b0100110000001011: data <= 8'b11111111;
		16'b0100110000001100: data <= 8'b11111111;
		16'b0100110000001101: data <= 8'b11111111;
		16'b0100110000001110: data <= 8'b11111111;
		16'b0100110000001111: data <= 8'b11111111;
		16'b0100110000010000: data <= 8'b11111111;
		16'b0100110000010001: data <= 8'b11111111;
		16'b0100110000010010: data <= 8'b11111111;
		16'b0100110000010011: data <= 8'b11111111;
		16'b0100110000010100: data <= 8'b11111111;
		16'b0100110000010101: data <= 8'b11111111;
		16'b0100110000010110: data <= 8'b11111111;
		16'b0100110000010111: data <= 8'b11111111;
		16'b0100110000011000: data <= 8'b11111111;
		16'b0100110000011001: data <= 8'b11111111;
		16'b0100110000011010: data <= 8'b11111111;
		16'b0100110000011011: data <= 8'b11111111;
		16'b0100110000011100: data <= 8'b11111111;
		16'b0100110000011101: data <= 8'b11111111;
		16'b0100110000011110: data <= 8'b11111111;
		16'b0100110000011111: data <= 8'b11111111;
		16'b0100110000100000: data <= 8'b11111111;
		16'b0100110000100001: data <= 8'b11111111;
		16'b0100110000100010: data <= 8'b11111111;
		16'b0100110000100011: data <= 8'b11111111;
		16'b0100110000100100: data <= 8'b11111111;
		16'b0100110000100101: data <= 8'b11111111;
		16'b0100110000100110: data <= 8'b11111111;
		16'b0100110000100111: data <= 8'b11111111;
		16'b0100110000101000: data <= 8'b11111111;
		16'b0100110000101001: data <= 8'b11111111;
		16'b0100110000101010: data <= 8'b11111111;
		16'b0100110000101011: data <= 8'b11111111;
		16'b0100110000101100: data <= 8'b11111111;
		16'b0100110000101101: data <= 8'b11111111;
		16'b0100110000101110: data <= 8'b11111111;
		16'b0100110000101111: data <= 8'b11111111;
		16'b0100110000110000: data <= 8'b11111111;
		16'b0100110000110001: data <= 8'b11111111;
		16'b0100110000110010: data <= 8'b11111111;
		16'b0100110000110011: data <= 8'b11111111;
		16'b0100110000110100: data <= 8'b11111111;
		16'b0100110000110101: data <= 8'b11111111;
		16'b0100110000110110: data <= 8'b11111111;
		16'b0100110000110111: data <= 8'b11111111;
		16'b0100110000111000: data <= 8'b11111111;
		16'b0100110000111001: data <= 8'b11111111;
		16'b0100110000111010: data <= 8'b11111111;
		16'b0100110000111011: data <= 8'b11111111;
		16'b0100110000111100: data <= 8'b11111111;
		16'b0100110000111101: data <= 8'b11111111;
		16'b0100110000111110: data <= 8'b11111111;
		16'b0100110000111111: data <= 8'b11111111;
		16'b0100110001000000: data <= 8'b11111111;
		16'b0100110001000001: data <= 8'b11111111;
		16'b0100110001000010: data <= 8'b11111111;
		16'b0100110001000011: data <= 8'b11111111;
		16'b0100110001000100: data <= 8'b11111111;
		16'b0100110001000101: data <= 8'b11111111;
		16'b0100110001000110: data <= 8'b11111111;
		16'b0100110001000111: data <= 8'b11111111;
		16'b0100110001001000: data <= 8'b11111111;
		16'b0100110001001001: data <= 8'b11111111;
		16'b0100110001001010: data <= 8'b11111111;
		16'b0100110001001011: data <= 8'b11111111;
		16'b0100110001001100: data <= 8'b11111111;
		16'b0100110001001101: data <= 8'b11111111;
		16'b0100110001001110: data <= 8'b11111111;
		16'b0100110001001111: data <= 8'b11111111;
		16'b0100110001010000: data <= 8'b11111111;
		16'b0100110001010001: data <= 8'b11111111;
		16'b0100110001010010: data <= 8'b11111111;
		16'b0100110001010011: data <= 8'b11111111;
		16'b0100110001010100: data <= 8'b11111111;
		16'b0100110001010101: data <= 8'b11111111;
		16'b0100110001010110: data <= 8'b11111111;
		16'b0100110001010111: data <= 8'b11111111;
		16'b0100110001011000: data <= 8'b11111111;
		16'b0100110001011001: data <= 8'b11111111;
		16'b0100110001011010: data <= 8'b11111111;
		16'b0100110001011011: data <= 8'b11111111;
		16'b0100110001011100: data <= 8'b11111111;
		16'b0100110001011101: data <= 8'b11111111;
		16'b0100110001011110: data <= 8'b11111111;
		16'b0100110001011111: data <= 8'b11111111;
		16'b0100110001100000: data <= 8'b11111111;
		16'b0100110001100001: data <= 8'b11111111;
		16'b0100110001100010: data <= 8'b11111111;
		16'b0100110001100011: data <= 8'b11111111;
		16'b0100110001100100: data <= 8'b11111111;
		16'b0100110001100101: data <= 8'b11111111;
		16'b0100110001100110: data <= 8'b11111111;
		16'b0100110001100111: data <= 8'b11111111;
		16'b0100110001101000: data <= 8'b11111111;
		16'b0100110001101001: data <= 8'b11111111;
		16'b0100110001101010: data <= 8'b11111111;
		16'b0100110001101011: data <= 8'b11111111;
		16'b0100110001101100: data <= 8'b11111111;
		16'b0100110001101101: data <= 8'b11111111;
		16'b0100110001101110: data <= 8'b11111111;
		16'b0100110001101111: data <= 8'b11111111;
		16'b0100110001110000: data <= 8'b11111111;
		16'b0100110001110001: data <= 8'b11111111;
		16'b0100110001110010: data <= 8'b11111111;
		16'b0100110001110011: data <= 8'b11111111;
		16'b0100110001110100: data <= 8'b11111111;
		16'b0100110001110101: data <= 8'b11111111;
		16'b0100110001110110: data <= 8'b11111111;
		16'b0100110001110111: data <= 8'b11111111;
		16'b0100110001111000: data <= 8'b11111111;
		16'b0100110001111001: data <= 8'b11111111;
		16'b0100110001111010: data <= 8'b11111111;
		16'b0100110001111011: data <= 8'b11111111;
		16'b0100110001111100: data <= 8'b11111111;
		16'b0100110001111101: data <= 8'b11111111;
		16'b0100110001111110: data <= 8'b11111111;
		16'b0100110001111111: data <= 8'b11111111;
		16'b0100110010000000: data <= 8'b11111111;
		16'b0100110010000001: data <= 8'b11111111;
		16'b0100110010000010: data <= 8'b11111111;
		16'b0100110010000011: data <= 8'b11111111;
		16'b0100110010000100: data <= 8'b11111111;
		16'b0100110010000101: data <= 8'b11111111;
		16'b0100110010000110: data <= 8'b11111111;
		16'b0100110010000111: data <= 8'b11111111;
		16'b0100110010001000: data <= 8'b11111111;
		16'b0100110010001001: data <= 8'b11111111;
		16'b0100110010001010: data <= 8'b11111111;
		16'b0100110010001011: data <= 8'b11111111;
		16'b0100110010001100: data <= 8'b11111111;
		16'b0100110010001101: data <= 8'b11111111;
		16'b0100110010001110: data <= 8'b11111111;
		16'b0100110010001111: data <= 8'b11111111;
		16'b0100110010010000: data <= 8'b11111111;
		16'b0100110010010001: data <= 8'b11111111;
		16'b0100110010010010: data <= 8'b11111111;
		16'b0100110010010011: data <= 8'b11111111;
		16'b0100110010010100: data <= 8'b11111111;
		16'b0100110010010101: data <= 8'b11111111;
		16'b0100110010010110: data <= 8'b11111111;
		16'b0100110010010111: data <= 8'b11111111;
		16'b0100110010011000: data <= 8'b11111111;
		16'b0100110010011001: data <= 8'b11111111;
		16'b0100110010011010: data <= 8'b11111111;
		16'b0100110010011011: data <= 8'b11111111;
		16'b0100110010011100: data <= 8'b11111111;
		16'b0100110010011101: data <= 8'b11111111;
		16'b0100110010011110: data <= 8'b11111111;
		16'b0100110010011111: data <= 8'b11111111;
		16'b0100110010100000: data <= 8'b11111111;
		16'b0100110010100001: data <= 8'b11111111;
		16'b0100110010100010: data <= 8'b11111111;
		16'b0100110010100011: data <= 8'b11111111;
		16'b0100110010100100: data <= 8'b11111111;
		16'b0100110010100101: data <= 8'b11111111;
		16'b0100110010100110: data <= 8'b11111111;
		16'b0100110010100111: data <= 8'b11111111;
		16'b0100110010101000: data <= 8'b11111111;
		16'b0100110010101001: data <= 8'b11111111;
		16'b0100110010101010: data <= 8'b11111111;
		16'b0100110010101011: data <= 8'b11111111;
		16'b0100110010101100: data <= 8'b11111111;
		16'b0100110010101101: data <= 8'b11111111;
		16'b0100110010101110: data <= 8'b11111111;
		16'b0100110010101111: data <= 8'b11111111;
		16'b0100110010110000: data <= 8'b11111111;
		16'b0100110010110001: data <= 8'b11111111;
		16'b0100110010110010: data <= 8'b11111111;
		16'b0100110010110011: data <= 8'b11111111;
		16'b0100110010110100: data <= 8'b11111111;
		16'b0100110010110101: data <= 8'b11111111;
		16'b0100110010110110: data <= 8'b11111111;
		16'b0100110010110111: data <= 8'b11111111;
		16'b0100110010111000: data <= 8'b11111111;
		16'b0100110010111001: data <= 8'b11111111;
		16'b0100110010111010: data <= 8'b11111111;
		16'b0100110010111011: data <= 8'b11111111;
		16'b0100110010111100: data <= 8'b11111111;
		16'b0100110010111101: data <= 8'b11111111;
		16'b0100110010111110: data <= 8'b11111111;
		16'b0100110010111111: data <= 8'b11111111;
		16'b0100110011000000: data <= 8'b11111111;
		16'b0100110011000001: data <= 8'b11111111;
		16'b0100110011000010: data <= 8'b11111111;
		16'b0100110011000011: data <= 8'b11111111;
		16'b0100110011000100: data <= 8'b11111111;
		16'b0100110011000101: data <= 8'b11111111;
		16'b0100110011000110: data <= 8'b11111111;
		16'b0100110011000111: data <= 8'b11111111;
		16'b0100110011001000: data <= 8'b11111111;
		16'b0100110011001001: data <= 8'b11111111;
		16'b0100110011001010: data <= 8'b11111111;
		16'b0100110011001011: data <= 8'b11111111;
		16'b0100110011001100: data <= 8'b11111111;
		16'b0100110011001101: data <= 8'b11111111;
		16'b0100110011001110: data <= 8'b11111111;
		16'b0100110011001111: data <= 8'b11111111;
		16'b0100110011010000: data <= 8'b11111111;
		16'b0100110011010001: data <= 8'b11111111;
		16'b0100110011010010: data <= 8'b11111111;
		16'b0100110011010011: data <= 8'b11111111;
		16'b0100110011010100: data <= 8'b11111111;
		16'b0100110011010101: data <= 8'b11111111;
		16'b0100110011010110: data <= 8'b11111111;
		16'b0100110011010111: data <= 8'b11111111;
		16'b0100110011011000: data <= 8'b11111111;
		16'b0100110011011001: data <= 8'b11111111;
		16'b0100110011011010: data <= 8'b11111111;
		16'b0100110011011011: data <= 8'b11111111;
		16'b0100110011011100: data <= 8'b11111111;
		16'b0100110011011101: data <= 8'b11111111;
		16'b0100110011011110: data <= 8'b11111111;
		16'b0100110011011111: data <= 8'b11111111;
		16'b0100110100101110: data <= 8'b11111111;
		16'b0100110100101111: data <= 8'b11111111;
		16'b0100110100110000: data <= 8'b11111111;
		16'b0100110100110001: data <= 8'b11111111;
		16'b0100110101111110: data <= 8'b11111111;
		16'b0100110101111111: data <= 8'b11111111;
		16'b0100110110000000: data <= 8'b11111111;
		16'b0100110110000001: data <= 8'b11111111;
		16'b0100111000011110: data <= 8'b11111111;
		16'b0100111000011111: data <= 8'b11111111;
		16'b0100111000100000: data <= 8'b11111111;
		16'b0100111000100001: data <= 8'b11111111;
		16'b0100111001101110: data <= 8'b11111111;
		16'b0100111001101111: data <= 8'b11111111;
		16'b0100111001110000: data <= 8'b11111111;
		16'b0100111001110001: data <= 8'b11111111;
		16'b0100111100001110: data <= 8'b11111111;
		16'b0100111100001111: data <= 8'b11111111;
		16'b0100111100010000: data <= 8'b11111111;
		16'b0100111100010001: data <= 8'b11111111;
		16'b0100111101011110: data <= 8'b11111111;
		16'b0100111101011111: data <= 8'b11111111;
		16'b0100111101100000: data <= 8'b11111111;
		16'b0100111101100001: data <= 8'b11111111;
		16'b0100111111111110: data <= 8'b11111111;
		16'b0100111111111111: data <= 8'b11111111;
		16'b0101000000000000: data <= 8'b11111111;
		16'b0101000000000001: data <= 8'b11111111;
		16'b0101000001001110: data <= 8'b11111111;
		16'b0101000001001111: data <= 8'b11111111;
		16'b0101000001010000: data <= 8'b11111111;
		16'b0101000001010001: data <= 8'b11111111;
		16'b0101000011101110: data <= 8'b11111111;
		16'b0101000011101111: data <= 8'b11111111;
		16'b0101000011110000: data <= 8'b11111111;
		16'b0101000011110001: data <= 8'b11111111;
		16'b0101000100111110: data <= 8'b11111111;
		16'b0101000100111111: data <= 8'b11111111;
		16'b0101000101000000: data <= 8'b11111111;
		16'b0101000101000001: data <= 8'b11111111;
		16'b0101000111011110: data <= 8'b11111111;
		16'b0101000111011111: data <= 8'b11111111;
		16'b0101000111100000: data <= 8'b11111111;
		16'b0101000111100001: data <= 8'b11111111;
		16'b0101001000101110: data <= 8'b11111111;
		16'b0101001000101111: data <= 8'b11111111;
		16'b0101001000110000: data <= 8'b11111111;
		16'b0101001000110001: data <= 8'b11111111;
		16'b0101001011001110: data <= 8'b11111111;
		16'b0101001011001111: data <= 8'b11111111;
		16'b0101001011010000: data <= 8'b11111111;
		16'b0101001011010001: data <= 8'b11111111;
		16'b0101001100011110: data <= 8'b11111111;
		16'b0101001100011111: data <= 8'b11111111;
		16'b0101001100100000: data <= 8'b11111111;
		16'b0101001100100001: data <= 8'b11111111;
		16'b0101001110111110: data <= 8'b11111111;
		16'b0101001110111111: data <= 8'b11111111;
		16'b0101001111000000: data <= 8'b11111111;
		16'b0101001111000001: data <= 8'b11111111;
		16'b0101010000001110: data <= 8'b11111111;
		16'b0101010000001111: data <= 8'b11111111;
		16'b0101010000010000: data <= 8'b11111111;
		16'b0101010000010001: data <= 8'b11111111;
		16'b0101010010101110: data <= 8'b11111111;
		16'b0101010010101111: data <= 8'b11111111;
		16'b0101010010110000: data <= 8'b11111111;
		16'b0101010010110001: data <= 8'b11111111;
		16'b0101010011111110: data <= 8'b11111111;
		16'b0101010011111111: data <= 8'b11111111;
		16'b0101010100000000: data <= 8'b11111111;
		16'b0101010100000001: data <= 8'b11111111;
		16'b0101010110011110: data <= 8'b11111111;
		16'b0101010110011111: data <= 8'b11111111;
		16'b0101010110100000: data <= 8'b11111111;
		16'b0101010110100001: data <= 8'b11111111;
		16'b0101010111101110: data <= 8'b11111111;
		16'b0101010111101111: data <= 8'b11111111;
		16'b0101010111110000: data <= 8'b11111111;
		16'b0101010111110001: data <= 8'b11111111;
		16'b0101011010001110: data <= 8'b11111111;
		16'b0101011010001111: data <= 8'b11111111;
		16'b0101011010010000: data <= 8'b11111111;
		16'b0101011010010001: data <= 8'b11111111;
		16'b0101011011011110: data <= 8'b11111111;
		16'b0101011011011111: data <= 8'b11111111;
		16'b0101011011100000: data <= 8'b11111111;
		16'b0101011011100001: data <= 8'b11111111;
		16'b0101011101111110: data <= 8'b11111111;
		16'b0101011101111111: data <= 8'b11111111;
		16'b0101011110000000: data <= 8'b11111111;
		16'b0101011110000001: data <= 8'b11111111;
		16'b0101011111001110: data <= 8'b11111111;
		16'b0101011111001111: data <= 8'b11111111;
		16'b0101011111010000: data <= 8'b11111111;
		16'b0101011111010001: data <= 8'b11111111;
		16'b0101100001101110: data <= 8'b11111111;
		16'b0101100001101111: data <= 8'b11111111;
		16'b0101100001110000: data <= 8'b11111111;
		16'b0101100001110001: data <= 8'b11111111;
		16'b0101100010111110: data <= 8'b11111111;
		16'b0101100010111111: data <= 8'b11111111;
		16'b0101100011000000: data <= 8'b11111111;
		16'b0101100011000001: data <= 8'b11111111;
		16'b0101100101011110: data <= 8'b11111111;
		16'b0101100101011111: data <= 8'b11111111;
		16'b0101100101100000: data <= 8'b11111111;
		16'b0101100101100001: data <= 8'b11111111;
		16'b0101100110101110: data <= 8'b11111111;
		16'b0101100110101111: data <= 8'b11111111;
		16'b0101100110110000: data <= 8'b11111111;
		16'b0101100110110001: data <= 8'b11111111;
		16'b0101101001001110: data <= 8'b11111111;
		16'b0101101001001111: data <= 8'b11111111;
		16'b0101101001010000: data <= 8'b11111111;
		16'b0101101001010001: data <= 8'b11111111;
		16'b0101101010011110: data <= 8'b11111111;
		16'b0101101010011111: data <= 8'b11111111;
		16'b0101101010100000: data <= 8'b11111111;
		16'b0101101010100001: data <= 8'b11111111;
		16'b0101101100111110: data <= 8'b11111111;
		16'b0101101100111111: data <= 8'b11111111;
		16'b0101101101000000: data <= 8'b11111111;
		16'b0101101101000001: data <= 8'b11111111;
		16'b0101101110001110: data <= 8'b11111111;
		16'b0101101110001111: data <= 8'b11111111;
		16'b0101101110010000: data <= 8'b11111111;
		16'b0101101110010001: data <= 8'b11111111;
		16'b0101110000101110: data <= 8'b11111111;
		16'b0101110000101111: data <= 8'b11111111;
		16'b0101110000110000: data <= 8'b11111111;
		16'b0101110000110001: data <= 8'b11111111;
		16'b0101110001111110: data <= 8'b11111111;
		16'b0101110001111111: data <= 8'b11111111;
		16'b0101110010000000: data <= 8'b11111111;
		16'b0101110010000001: data <= 8'b11111111;
		16'b0101110100011110: data <= 8'b11111111;
		16'b0101110100011111: data <= 8'b11111111;
		16'b0101110100100000: data <= 8'b11111111;
		16'b0101110100100001: data <= 8'b11111111;
		16'b0101110101101110: data <= 8'b11111111;
		16'b0101110101101111: data <= 8'b11111111;
		16'b0101110101110000: data <= 8'b11111111;
		16'b0101110101110001: data <= 8'b11111111;
		16'b0101111000001110: data <= 8'b11111111;
		16'b0101111000001111: data <= 8'b11111111;
		16'b0101111000010000: data <= 8'b11111111;
		16'b0101111000010001: data <= 8'b11111111;
		16'b0101111001011110: data <= 8'b11111111;
		16'b0101111001011111: data <= 8'b11111111;
		16'b0101111001100000: data <= 8'b11111111;
		16'b0101111001100001: data <= 8'b11111111;
		16'b0101111011111110: data <= 8'b11111111;
		16'b0101111011111111: data <= 8'b11111111;
		16'b0101111100000000: data <= 8'b11111111;
		16'b0101111100000001: data <= 8'b11111111;
		16'b0101111101001110: data <= 8'b11111111;
		16'b0101111101001111: data <= 8'b11111111;
		16'b0101111101010000: data <= 8'b11111111;
		16'b0101111101010001: data <= 8'b11111111;
		16'b0101111111101110: data <= 8'b11111111;
		16'b0101111111101111: data <= 8'b11111111;
		16'b0101111111110000: data <= 8'b11111111;
		16'b0101111111110001: data <= 8'b11111111;
		16'b0110000000111110: data <= 8'b11111111;
		16'b0110000000111111: data <= 8'b11111111;
		16'b0110000001000000: data <= 8'b11111111;
		16'b0110000001000001: data <= 8'b11111111;
		16'b0110000011011110: data <= 8'b11111111;
		16'b0110000011011111: data <= 8'b11111111;
		16'b0110000011100000: data <= 8'b11111111;
		16'b0110000011100001: data <= 8'b11111111;
		16'b0110000100101110: data <= 8'b11111111;
		16'b0110000100101111: data <= 8'b11111111;
		16'b0110000100110000: data <= 8'b11111111;
		16'b0110000100110001: data <= 8'b11111111;
		16'b0110000111001110: data <= 8'b11111111;
		16'b0110000111001111: data <= 8'b11111111;
		16'b0110000111010000: data <= 8'b11111111;
		16'b0110000111010001: data <= 8'b11111111;
		16'b0110001000011110: data <= 8'b11111111;
		16'b0110001000011111: data <= 8'b11111111;
		16'b0110001000100000: data <= 8'b11111111;
		16'b0110001000100001: data <= 8'b11111111;
		16'b0110001010111110: data <= 8'b11111111;
		16'b0110001010111111: data <= 8'b11111111;
		16'b0110001011000000: data <= 8'b11111111;
		16'b0110001011000001: data <= 8'b11111111;
		16'b0110001100001110: data <= 8'b11111111;
		16'b0110001100001111: data <= 8'b11111111;
		16'b0110001100010000: data <= 8'b11111111;
		16'b0110001100010001: data <= 8'b11111111;
		16'b0110001110101110: data <= 8'b11111111;
		16'b0110001110101111: data <= 8'b11111111;
		16'b0110001110110000: data <= 8'b11111111;
		16'b0110001110110001: data <= 8'b11111111;
		16'b0110001111111110: data <= 8'b11111111;
		16'b0110001111111111: data <= 8'b11111111;
		16'b0110010000000000: data <= 8'b11111111;
		16'b0110010000000001: data <= 8'b11111111;
		16'b0110010010011110: data <= 8'b11111111;
		16'b0110010010011111: data <= 8'b11111111;
		16'b0110010010100000: data <= 8'b11111111;
		16'b0110010010100001: data <= 8'b11111111;
		16'b0110010011101110: data <= 8'b11111111;
		16'b0110010011101111: data <= 8'b11111111;
		16'b0110010011110000: data <= 8'b11111111;
		16'b0110010011110001: data <= 8'b11111111;
		16'b0110010110001110: data <= 8'b11111111;
		16'b0110010110001111: data <= 8'b11111111;
		16'b0110010110010000: data <= 8'b11111111;
		16'b0110010110010001: data <= 8'b11111111;
		16'b0110010111011110: data <= 8'b11111111;
		16'b0110010111011111: data <= 8'b11111111;
		16'b0110010111100000: data <= 8'b11111111;
		16'b0110010111100001: data <= 8'b11111111;
		16'b0110011001111110: data <= 8'b11111111;
		16'b0110011001111111: data <= 8'b11111111;
		16'b0110011010000000: data <= 8'b11111111;
		16'b0110011010000001: data <= 8'b11111111;
		16'b0110011011001110: data <= 8'b11111111;
		16'b0110011011001111: data <= 8'b11111111;
		16'b0110011011010000: data <= 8'b11111111;
		16'b0110011011010001: data <= 8'b11111111;
		16'b0110011101101110: data <= 8'b11111111;
		16'b0110011101101111: data <= 8'b11111111;
		16'b0110011101110000: data <= 8'b11111111;
		16'b0110011101110001: data <= 8'b11111111;
		16'b0110011110111110: data <= 8'b11111111;
		16'b0110011110111111: data <= 8'b11111111;
		16'b0110011111000000: data <= 8'b11111111;
		16'b0110011111000001: data <= 8'b11111111;
		16'b0110100001011110: data <= 8'b11111111;
		16'b0110100001011111: data <= 8'b11111111;
		16'b0110100001100000: data <= 8'b11111111;
		16'b0110100001100001: data <= 8'b11111111;
		16'b0110100010101110: data <= 8'b11111111;
		16'b0110100010101111: data <= 8'b11111111;
		16'b0110100010110000: data <= 8'b11111111;
		16'b0110100010110001: data <= 8'b11111111;
		16'b0110100101001110: data <= 8'b11111111;
		16'b0110100101001111: data <= 8'b11111111;
		16'b0110100101010000: data <= 8'b11111111;
		16'b0110100101010001: data <= 8'b11111111;
		16'b0110100110011110: data <= 8'b11111111;
		16'b0110100110011111: data <= 8'b11111111;
		16'b0110100110100000: data <= 8'b11111111;
		16'b0110100110100001: data <= 8'b11111111;
		16'b0110101000111110: data <= 8'b11111111;
		16'b0110101000111111: data <= 8'b11111111;
		16'b0110101001000000: data <= 8'b11111111;
		16'b0110101001000001: data <= 8'b11111111;
		16'b0110101010001110: data <= 8'b11111111;
		16'b0110101010001111: data <= 8'b11111111;
		16'b0110101010010000: data <= 8'b11111111;
		16'b0110101010010001: data <= 8'b11111111;
		16'b0110101100101110: data <= 8'b11111111;
		16'b0110101100101111: data <= 8'b11111111;
		16'b0110101100110000: data <= 8'b11111111;
		16'b0110101100110001: data <= 8'b11111111;
		16'b0110101101111110: data <= 8'b11111111;
		16'b0110101101111111: data <= 8'b11111111;
		16'b0110101110000000: data <= 8'b11111111;
		16'b0110101110000001: data <= 8'b11111111;
		16'b0110110000011110: data <= 8'b11111111;
		16'b0110110000011111: data <= 8'b11111111;
		16'b0110110000100000: data <= 8'b11111111;
		16'b0110110000100001: data <= 8'b11111111;
		16'b0110110001101110: data <= 8'b11111111;
		16'b0110110001101111: data <= 8'b11111111;
		16'b0110110001110000: data <= 8'b11111111;
		16'b0110110001110001: data <= 8'b11111111;
		16'b0110110100001110: data <= 8'b11111111;
		16'b0110110100001111: data <= 8'b11111111;
		16'b0110110100010000: data <= 8'b11111111;
		16'b0110110100010001: data <= 8'b11111111;
		16'b0110110101011110: data <= 8'b11111111;
		16'b0110110101011111: data <= 8'b11111111;
		16'b0110110101100000: data <= 8'b11111111;
		16'b0110110101100001: data <= 8'b11111111;
		16'b0110110111111110: data <= 8'b11111111;
		16'b0110110111111111: data <= 8'b11111111;
		16'b0110111000000000: data <= 8'b11111111;
		16'b0110111000000001: data <= 8'b11111111;
		16'b0110111001001110: data <= 8'b11111111;
		16'b0110111001001111: data <= 8'b11111111;
		16'b0110111001010000: data <= 8'b11111111;
		16'b0110111001010001: data <= 8'b11111111;
		16'b0110111011101110: data <= 8'b11111111;
		16'b0110111011101111: data <= 8'b11111111;
		16'b0110111011110000: data <= 8'b11111111;
		16'b0110111011110001: data <= 8'b11111111;
		16'b0110111100111110: data <= 8'b11111111;
		16'b0110111100111111: data <= 8'b11111111;
		16'b0110111101000000: data <= 8'b11111111;
		16'b0110111101000001: data <= 8'b11111111;
		16'b0110111111011110: data <= 8'b11111111;
		16'b0110111111011111: data <= 8'b11111111;
		16'b0110111111100000: data <= 8'b11111111;
		16'b0110111111100001: data <= 8'b11111111;
		16'b0111000000101110: data <= 8'b11111111;
		16'b0111000000101111: data <= 8'b11111111;
		16'b0111000000110000: data <= 8'b11111111;
		16'b0111000000110001: data <= 8'b11111111;
		16'b0111000011001110: data <= 8'b11111111;
		16'b0111000011001111: data <= 8'b11111111;
		16'b0111000011010000: data <= 8'b11111111;
		16'b0111000011010001: data <= 8'b11111111;
		16'b0111000100011110: data <= 8'b11111111;
		16'b0111000100011111: data <= 8'b11111111;
		16'b0111000100100000: data <= 8'b11111111;
		16'b0111000100100001: data <= 8'b11111111;
		16'b0111000110111110: data <= 8'b11111111;
		16'b0111000110111111: data <= 8'b11111111;
		16'b0111000111000000: data <= 8'b11111111;
		16'b0111000111000001: data <= 8'b11111111;
		16'b0111001000001110: data <= 8'b11111111;
		16'b0111001000001111: data <= 8'b11111111;
		16'b0111001000010000: data <= 8'b11111111;
		16'b0111001000010001: data <= 8'b11111111;
		16'b0111001010101110: data <= 8'b11111111;
		16'b0111001010101111: data <= 8'b11111111;
		16'b0111001010110000: data <= 8'b11111111;
		16'b0111001010110001: data <= 8'b11111111;
		16'b0111001011111110: data <= 8'b11111111;
		16'b0111001011111111: data <= 8'b11111111;
		16'b0111001100000000: data <= 8'b11111111;
		16'b0111001100000001: data <= 8'b11111111;
		16'b0111001110011110: data <= 8'b11111111;
		16'b0111001110011111: data <= 8'b11111111;
		16'b0111001110100000: data <= 8'b11111111;
		16'b0111001110100001: data <= 8'b11111111;
		16'b0111001111101110: data <= 8'b11111111;
		16'b0111001111101111: data <= 8'b11111111;
		16'b0111001111110000: data <= 8'b11111111;
		16'b0111001111110001: data <= 8'b11111111;
		16'b0111010010001110: data <= 8'b11111111;
		16'b0111010010001111: data <= 8'b11111111;
		16'b0111010010010000: data <= 8'b11111111;
		16'b0111010010010001: data <= 8'b11111111;
		16'b0111010011011110: data <= 8'b11111111;
		16'b0111010011011111: data <= 8'b11111111;
		16'b0111010011100000: data <= 8'b11111111;
		16'b0111010011100001: data <= 8'b11111111;
		16'b0111010101111110: data <= 8'b11111111;
		16'b0111010101111111: data <= 8'b11111111;
		16'b0111010110000000: data <= 8'b11111111;
		16'b0111010110000001: data <= 8'b11111111;
		16'b0111010111001110: data <= 8'b11111111;
		16'b0111010111001111: data <= 8'b11111111;
		16'b0111010111010000: data <= 8'b11111111;
		16'b0111010111010001: data <= 8'b11111111;
		16'b0111011001101110: data <= 8'b11111111;
		16'b0111011001101111: data <= 8'b11111111;
		16'b0111011001110000: data <= 8'b11111111;
		16'b0111011001110001: data <= 8'b11111111;
		16'b0111011010111110: data <= 8'b11111111;
		16'b0111011010111111: data <= 8'b11111111;
		16'b0111011011000000: data <= 8'b11111111;
		16'b0111011011000001: data <= 8'b11111111;
		16'b0111011101011110: data <= 8'b11111111;
		16'b0111011101011111: data <= 8'b11111111;
		16'b0111011101100000: data <= 8'b11111111;
		16'b0111011101100001: data <= 8'b11111111;
		16'b0111011110101110: data <= 8'b11111111;
		16'b0111011110101111: data <= 8'b11111111;
		16'b0111011110110000: data <= 8'b11111111;
		16'b0111011110110001: data <= 8'b11111111;
		16'b0111100001001110: data <= 8'b11111111;
		16'b0111100001001111: data <= 8'b11111111;
		16'b0111100001010000: data <= 8'b11111111;
		16'b0111100001010001: data <= 8'b11111111;
		16'b0111100010011110: data <= 8'b11111111;
		16'b0111100010011111: data <= 8'b11111111;
		16'b0111100010100000: data <= 8'b11111111;
		16'b0111100010100001: data <= 8'b11111111;
		16'b0111100100111110: data <= 8'b11111111;
		16'b0111100100111111: data <= 8'b11111111;
		16'b0111100101000000: data <= 8'b11111111;
		16'b0111100101000001: data <= 8'b11111111;
		16'b0111100110001110: data <= 8'b11111111;
		16'b0111100110001111: data <= 8'b11111111;
		16'b0111100110010000: data <= 8'b11111111;
		16'b0111100110010001: data <= 8'b11111111;
		16'b0111101000101110: data <= 8'b11111111;
		16'b0111101000101111: data <= 8'b11111111;
		16'b0111101000110000: data <= 8'b11111111;
		16'b0111101000110001: data <= 8'b11111111;
		16'b0111101001111110: data <= 8'b11111111;
		16'b0111101001111111: data <= 8'b11111111;
		16'b0111101010000000: data <= 8'b11111111;
		16'b0111101010000001: data <= 8'b11111111;
		16'b0111101100011110: data <= 8'b11111111;
		16'b0111101100011111: data <= 8'b11111111;
		16'b0111101100100000: data <= 8'b11111111;
		16'b0111101100100001: data <= 8'b11111111;
		16'b0111101101101110: data <= 8'b11111111;
		16'b0111101101101111: data <= 8'b11111111;
		16'b0111101101110000: data <= 8'b11111111;
		16'b0111101101110001: data <= 8'b11111111;
		16'b0111110000001110: data <= 8'b11111111;
		16'b0111110000001111: data <= 8'b11111111;
		16'b0111110000010000: data <= 8'b11111111;
		16'b0111110000010001: data <= 8'b11111111;
		16'b0111110001011110: data <= 8'b11111111;
		16'b0111110001011111: data <= 8'b11111111;
		16'b0111110001100000: data <= 8'b11111111;
		16'b0111110001100001: data <= 8'b11111111;
		16'b0111110011111110: data <= 8'b11111111;
		16'b0111110011111111: data <= 8'b11111111;
		16'b0111110100000000: data <= 8'b11111111;
		16'b0111110100000001: data <= 8'b11111111;
		16'b0111110101001110: data <= 8'b11111111;
		16'b0111110101001111: data <= 8'b11111111;
		16'b0111110101010000: data <= 8'b11111111;
		16'b0111110101010001: data <= 8'b11111111;
		16'b0111110111101110: data <= 8'b11111111;
		16'b0111110111101111: data <= 8'b11111111;
		16'b0111110111110000: data <= 8'b11111111;
		16'b0111110111110001: data <= 8'b11111111;
		16'b0111111000111110: data <= 8'b11111111;
		16'b0111111000111111: data <= 8'b11111111;
		16'b0111111001000000: data <= 8'b11111111;
		16'b0111111001000001: data <= 8'b11111111;
		16'b0111111011011110: data <= 8'b11111111;
		16'b0111111011011111: data <= 8'b11111111;
		16'b0111111011100000: data <= 8'b11111111;
		16'b0111111011100001: data <= 8'b11111111;
		16'b0111111100101110: data <= 8'b11111111;
		16'b0111111100101111: data <= 8'b11111111;
		16'b0111111100110000: data <= 8'b11111111;
		16'b0111111100110001: data <= 8'b11111111;
		16'b0111111111001110: data <= 8'b11111111;
		16'b0111111111001111: data <= 8'b11111111;
		16'b0111111111010000: data <= 8'b11111111;
		16'b0111111111010001: data <= 8'b11111111;
		16'b1000000000011110: data <= 8'b11111111;
		16'b1000000000011111: data <= 8'b11111111;
		16'b1000000000100000: data <= 8'b11111111;
		16'b1000000000100001: data <= 8'b11111111;
		16'b1000000010111110: data <= 8'b11111111;
		16'b1000000010111111: data <= 8'b11111111;
		16'b1000000011000000: data <= 8'b11111111;
		16'b1000000011000001: data <= 8'b11111111;
		16'b1000000100001110: data <= 8'b11111111;
		16'b1000000100001111: data <= 8'b11111111;
		16'b1000000100010000: data <= 8'b11111111;
		16'b1000000100010001: data <= 8'b11111111;
		16'b1000000110101110: data <= 8'b11111111;
		16'b1000000110101111: data <= 8'b11111111;
		16'b1000000110110000: data <= 8'b11111111;
		16'b1000000110110001: data <= 8'b11111111;
		16'b1000000111111110: data <= 8'b11111111;
		16'b1000000111111111: data <= 8'b11111111;
		16'b1000001000000000: data <= 8'b11111111;
		16'b1000001000000001: data <= 8'b11111111;
		16'b1000001010011110: data <= 8'b11111111;
		16'b1000001010011111: data <= 8'b11111111;
		16'b1000001010100000: data <= 8'b11111111;
		16'b1000001010100001: data <= 8'b11111111;
		16'b1000001011101110: data <= 8'b11111111;
		16'b1000001011101111: data <= 8'b11111111;
		16'b1000001011110000: data <= 8'b11111111;
		16'b1000001011110001: data <= 8'b11111111;
		16'b1000001110001110: data <= 8'b11111111;
		16'b1000001110001111: data <= 8'b11111111;
		16'b1000001110010000: data <= 8'b11111111;
		16'b1000001110010001: data <= 8'b11111111;
		16'b1000001111011110: data <= 8'b11111111;
		16'b1000001111011111: data <= 8'b11111111;
		16'b1000001111100000: data <= 8'b11111111;
		16'b1000001111100001: data <= 8'b11111111;
		16'b1000010001111110: data <= 8'b11111111;
		16'b1000010001111111: data <= 8'b11111111;
		16'b1000010010000000: data <= 8'b11111111;
		16'b1000010010000001: data <= 8'b11111111;
		16'b1000010011001110: data <= 8'b11111111;
		16'b1000010011001111: data <= 8'b11111111;
		16'b1000010011010000: data <= 8'b11111111;
		16'b1000010011010001: data <= 8'b11111111;
		16'b1000010101101110: data <= 8'b11111111;
		16'b1000010101101111: data <= 8'b11111111;
		16'b1000010101110000: data <= 8'b11111111;
		16'b1000010101110001: data <= 8'b11111111;
		16'b1000010110111110: data <= 8'b11111111;
		16'b1000010110111111: data <= 8'b11111111;
		16'b1000010111000000: data <= 8'b11111111;
		16'b1000010111000001: data <= 8'b11111111;
		16'b1000011001011110: data <= 8'b11111111;
		16'b1000011001011111: data <= 8'b11111111;
		16'b1000011001100000: data <= 8'b11111111;
		16'b1000011001100001: data <= 8'b11111111;
		16'b1000011010101110: data <= 8'b11111111;
		16'b1000011010101111: data <= 8'b11111111;
		16'b1000011010110000: data <= 8'b11111111;
		16'b1000011010110001: data <= 8'b11111111;
		16'b1000011101001110: data <= 8'b11111111;
		16'b1000011101001111: data <= 8'b11111111;
		16'b1000011101010000: data <= 8'b11111111;
		16'b1000011101010001: data <= 8'b11111111;
		16'b1000011110011110: data <= 8'b11111111;
		16'b1000011110011111: data <= 8'b11111111;
		16'b1000011110100000: data <= 8'b11111111;
		16'b1000011110100001: data <= 8'b11111111;
		16'b1000100000111110: data <= 8'b11111111;
		16'b1000100000111111: data <= 8'b11111111;
		16'b1000100001000000: data <= 8'b11111111;
		16'b1000100001000001: data <= 8'b11111111;
		16'b1000100010001110: data <= 8'b11111111;
		16'b1000100010001111: data <= 8'b11111111;
		16'b1000100010010000: data <= 8'b11111111;
		16'b1000100010010001: data <= 8'b11111111;
		16'b1000100100101110: data <= 8'b11111111;
		16'b1000100100101111: data <= 8'b11111111;
		16'b1000100100110000: data <= 8'b11111111;
		16'b1000100100110001: data <= 8'b11111111;
		16'b1000100101111110: data <= 8'b11111111;
		16'b1000100101111111: data <= 8'b11111111;
		16'b1000100110000000: data <= 8'b11111111;
		16'b1000100110000001: data <= 8'b11111111;
		16'b1000101000011110: data <= 8'b11111111;
		16'b1000101000011111: data <= 8'b11111111;
		16'b1000101000100000: data <= 8'b11111111;
		16'b1000101000100001: data <= 8'b11111111;
		16'b1000101001101110: data <= 8'b11111111;
		16'b1000101001101111: data <= 8'b11111111;
		16'b1000101001110000: data <= 8'b11111111;
		16'b1000101001110001: data <= 8'b11111111;
		16'b1000101100001110: data <= 8'b11111111;
		16'b1000101100001111: data <= 8'b11111111;
		16'b1000101100010000: data <= 8'b11111111;
		16'b1000101100010001: data <= 8'b11111111;
		16'b1000101101011110: data <= 8'b11111111;
		16'b1000101101011111: data <= 8'b11111111;
		16'b1000101101100000: data <= 8'b11111111;
		16'b1000101101100001: data <= 8'b11111111;
		16'b1000101111111110: data <= 8'b11111111;
		16'b1000101111111111: data <= 8'b11111111;
		16'b1000110000000000: data <= 8'b11111111;
		16'b1000110000000001: data <= 8'b11111111;
		16'b1000110001001110: data <= 8'b11111111;
		16'b1000110001001111: data <= 8'b11111111;
		16'b1000110001010000: data <= 8'b11111111;
		16'b1000110001010001: data <= 8'b11111111;
		16'b1000110011101110: data <= 8'b11111111;
		16'b1000110011101111: data <= 8'b11111111;
		16'b1000110011110000: data <= 8'b11111111;
		16'b1000110011110001: data <= 8'b11111111;
		16'b1000110100111110: data <= 8'b11111111;
		16'b1000110100111111: data <= 8'b11111111;
		16'b1000110101000000: data <= 8'b11111111;
		16'b1000110101000001: data <= 8'b11111111;
		16'b1000110111011110: data <= 8'b11111111;
		16'b1000110111011111: data <= 8'b11111111;
		16'b1000110111100000: data <= 8'b11111111;
		16'b1000110111100001: data <= 8'b11111111;
		16'b1000111000101110: data <= 8'b11111111;
		16'b1000111000101111: data <= 8'b11111111;
		16'b1000111000110000: data <= 8'b11111111;
		16'b1000111000110001: data <= 8'b11111111;
		16'b1000111011001110: data <= 8'b11111111;
		16'b1000111011001111: data <= 8'b11111111;
		16'b1000111011010000: data <= 8'b11111111;
		16'b1000111011010001: data <= 8'b11111111;
		16'b1000111100011110: data <= 8'b11111111;
		16'b1000111100011111: data <= 8'b11111111;
		16'b1000111100100000: data <= 8'b11111111;
		16'b1000111100100001: data <= 8'b11111111;
		16'b1000111110111110: data <= 8'b11111111;
		16'b1000111110111111: data <= 8'b11111111;
		16'b1000111111000000: data <= 8'b11111111;
		16'b1000111111000001: data <= 8'b11111111;
		16'b1001000000001110: data <= 8'b11111111;
		16'b1001000000001111: data <= 8'b11111111;
		16'b1001000000010000: data <= 8'b11111111;
		16'b1001000000010001: data <= 8'b11111111;
		16'b1001000010101110: data <= 8'b11111111;
		16'b1001000010101111: data <= 8'b11111111;
		16'b1001000010110000: data <= 8'b11111111;
		16'b1001000010110001: data <= 8'b11111111;
		16'b1001000011111110: data <= 8'b11111111;
		16'b1001000011111111: data <= 8'b11111111;
		16'b1001000100000000: data <= 8'b11111111;
		16'b1001000100000001: data <= 8'b11111111;
		16'b1001000110011110: data <= 8'b11111111;
		16'b1001000110011111: data <= 8'b11111111;
		16'b1001000110100000: data <= 8'b11111111;
		16'b1001000110100001: data <= 8'b11111111;
		16'b1001000111101110: data <= 8'b11111111;
		16'b1001000111101111: data <= 8'b11111111;
		16'b1001000111110000: data <= 8'b11111111;
		16'b1001000111110001: data <= 8'b11111111;
		16'b1001001010001110: data <= 8'b11111111;
		16'b1001001010001111: data <= 8'b11111111;
		16'b1001001010010000: data <= 8'b11111111;
		16'b1001001010010001: data <= 8'b11111111;
		16'b1001001011011110: data <= 8'b11111111;
		16'b1001001011011111: data <= 8'b11111111;
		16'b1001001011100000: data <= 8'b11111111;
		16'b1001001011100001: data <= 8'b11111111;
		16'b1001001101111110: data <= 8'b11111111;
		16'b1001001101111111: data <= 8'b11111111;
		16'b1001001110000000: data <= 8'b11111111;
		16'b1001001110000001: data <= 8'b11111111;
		16'b1001001111001110: data <= 8'b11111111;
		16'b1001001111001111: data <= 8'b11111111;
		16'b1001001111010000: data <= 8'b11111111;
		16'b1001001111010001: data <= 8'b11111111;
		16'b1001010000100000: data <= 8'b11111111;
		16'b1001010000100001: data <= 8'b11111111;
		16'b1001010000100010: data <= 8'b11111111;
		16'b1001010000100011: data <= 8'b11111111;
		16'b1001010000100100: data <= 8'b11111111;
		16'b1001010000100101: data <= 8'b11111111;
		16'b1001010000100110: data <= 8'b11111111;
		16'b1001010000100111: data <= 8'b11111111;
		16'b1001010000101000: data <= 8'b11111111;
		16'b1001010000101001: data <= 8'b11111111;
		16'b1001010000101010: data <= 8'b11111111;
		16'b1001010000101011: data <= 8'b11111111;
		16'b1001010000101100: data <= 8'b11111111;
		16'b1001010000101101: data <= 8'b11111111;
		16'b1001010000101110: data <= 8'b11111111;
		16'b1001010000101111: data <= 8'b11111111;
		16'b1001010000110000: data <= 8'b11111111;
		16'b1001010000110001: data <= 8'b11111111;
		16'b1001010000110010: data <= 8'b11111111;
		16'b1001010000110011: data <= 8'b11111111;
		16'b1001010000110100: data <= 8'b11111111;
		16'b1001010000110101: data <= 8'b11111111;
		16'b1001010000110110: data <= 8'b11111111;
		16'b1001010000110111: data <= 8'b11111111;
		16'b1001010000111000: data <= 8'b11111111;
		16'b1001010000111001: data <= 8'b11111111;
		16'b1001010000111010: data <= 8'b11111111;
		16'b1001010000111011: data <= 8'b11111111;
		16'b1001010000111100: data <= 8'b11111111;
		16'b1001010000111101: data <= 8'b11111111;
		16'b1001010000111110: data <= 8'b11111111;
		16'b1001010000111111: data <= 8'b11111111;
		16'b1001010001000000: data <= 8'b11111111;
		16'b1001010001000001: data <= 8'b11111111;
		16'b1001010001000010: data <= 8'b11111111;
		16'b1001010001000011: data <= 8'b11111111;
		16'b1001010001000100: data <= 8'b11111111;
		16'b1001010001000101: data <= 8'b11111111;
		16'b1001010001000110: data <= 8'b11111111;
		16'b1001010001000111: data <= 8'b11111111;
		16'b1001010001001000: data <= 8'b11111111;
		16'b1001010001001001: data <= 8'b11111111;
		16'b1001010001001010: data <= 8'b11111111;
		16'b1001010001001011: data <= 8'b11111111;
		16'b1001010001001100: data <= 8'b11111111;
		16'b1001010001001101: data <= 8'b11111111;
		16'b1001010001001110: data <= 8'b11111111;
		16'b1001010001001111: data <= 8'b11111111;
		16'b1001010001010000: data <= 8'b11111111;
		16'b1001010001010001: data <= 8'b11111111;
		16'b1001010001010010: data <= 8'b11111111;
		16'b1001010001010011: data <= 8'b11111111;
		16'b1001010001010100: data <= 8'b11111111;
		16'b1001010001010101: data <= 8'b11111111;
		16'b1001010001010110: data <= 8'b11111111;
		16'b1001010001010111: data <= 8'b11111111;
		16'b1001010001011000: data <= 8'b11111111;
		16'b1001010001011001: data <= 8'b11111111;
		16'b1001010001011010: data <= 8'b11111111;
		16'b1001010001011011: data <= 8'b11111111;
		16'b1001010001011100: data <= 8'b11111111;
		16'b1001010001011101: data <= 8'b11111111;
		16'b1001010001011110: data <= 8'b11111111;
		16'b1001010001011111: data <= 8'b11111111;
		16'b1001010001100000: data <= 8'b11111111;
		16'b1001010001100001: data <= 8'b11111111;
		16'b1001010001100010: data <= 8'b11111111;
		16'b1001010001100011: data <= 8'b11111111;
		16'b1001010001100100: data <= 8'b11111111;
		16'b1001010001100101: data <= 8'b11111111;
		16'b1001010001100110: data <= 8'b11111111;
		16'b1001010001100111: data <= 8'b11111111;
		16'b1001010001101000: data <= 8'b11111111;
		16'b1001010001101001: data <= 8'b11111111;
		16'b1001010001101010: data <= 8'b11111111;
		16'b1001010001101011: data <= 8'b11111111;
		16'b1001010001101100: data <= 8'b11111111;
		16'b1001010001101101: data <= 8'b11111111;
		16'b1001010001101110: data <= 8'b11111111;
		16'b1001010001101111: data <= 8'b11111111;
		16'b1001010001110000: data <= 8'b11111111;
		16'b1001010001110001: data <= 8'b11111111;
		16'b1001010001110010: data <= 8'b11111111;
		16'b1001010001110011: data <= 8'b11111111;
		16'b1001010001110100: data <= 8'b11111111;
		16'b1001010001110101: data <= 8'b11111111;
		16'b1001010001110110: data <= 8'b11111111;
		16'b1001010001110111: data <= 8'b11111111;
		16'b1001010001111000: data <= 8'b11111111;
		16'b1001010001111001: data <= 8'b11111111;
		16'b1001010001111010: data <= 8'b11111111;
		16'b1001010001111011: data <= 8'b11111111;
		16'b1001010001111100: data <= 8'b11111111;
		16'b1001010001111101: data <= 8'b11111111;
		16'b1001010001111110: data <= 8'b11111111;
		16'b1001010001111111: data <= 8'b11111111;
		16'b1001010010000000: data <= 8'b11111111;
		16'b1001010010000001: data <= 8'b11111111;
		16'b1001010010000010: data <= 8'b11111111;
		16'b1001010010000011: data <= 8'b11111111;
		16'b1001010010000100: data <= 8'b11111111;
		16'b1001010010000101: data <= 8'b11111111;
		16'b1001010010000110: data <= 8'b11111111;
		16'b1001010010000111: data <= 8'b11111111;
		16'b1001010010001000: data <= 8'b11111111;
		16'b1001010010001001: data <= 8'b11111111;
		16'b1001010010001010: data <= 8'b11111111;
		16'b1001010010001011: data <= 8'b11111111;
		16'b1001010010001100: data <= 8'b11111111;
		16'b1001010010001101: data <= 8'b11111111;
		16'b1001010010001110: data <= 8'b11111111;
		16'b1001010010001111: data <= 8'b11111111;
		16'b1001010010010000: data <= 8'b11111111;
		16'b1001010010010001: data <= 8'b11111111;
		16'b1001010010010010: data <= 8'b11111111;
		16'b1001010010010011: data <= 8'b11111111;
		16'b1001010010010100: data <= 8'b11111111;
		16'b1001010010010101: data <= 8'b11111111;
		16'b1001010010010110: data <= 8'b11111111;
		16'b1001010010010111: data <= 8'b11111111;
		16'b1001010010011000: data <= 8'b11111111;
		16'b1001010010011001: data <= 8'b11111111;
		16'b1001010010011010: data <= 8'b11111111;
		16'b1001010010011011: data <= 8'b11111111;
		16'b1001010010011100: data <= 8'b11111111;
		16'b1001010010011101: data <= 8'b11111111;
		16'b1001010010011110: data <= 8'b11111111;
		16'b1001010010011111: data <= 8'b11111111;
		16'b1001010010100000: data <= 8'b11111111;
		16'b1001010010100001: data <= 8'b11111111;
		16'b1001010010100010: data <= 8'b11111111;
		16'b1001010010100011: data <= 8'b11111111;
		16'b1001010010100100: data <= 8'b11111111;
		16'b1001010010100101: data <= 8'b11111111;
		16'b1001010010100110: data <= 8'b11111111;
		16'b1001010010100111: data <= 8'b11111111;
		16'b1001010010101000: data <= 8'b11111111;
		16'b1001010010101001: data <= 8'b11111111;
		16'b1001010010101010: data <= 8'b11111111;
		16'b1001010010101011: data <= 8'b11111111;
		16'b1001010010101100: data <= 8'b11111111;
		16'b1001010010101101: data <= 8'b11111111;
		16'b1001010010101110: data <= 8'b11111111;
		16'b1001010010101111: data <= 8'b11111111;
		16'b1001010010110000: data <= 8'b11111111;
		16'b1001010010110001: data <= 8'b11111111;
		16'b1001010010110010: data <= 8'b11111111;
		16'b1001010010110011: data <= 8'b11111111;
		16'b1001010010110100: data <= 8'b11111111;
		16'b1001010010110101: data <= 8'b11111111;
		16'b1001010010110110: data <= 8'b11111111;
		16'b1001010010110111: data <= 8'b11111111;
		16'b1001010010111000: data <= 8'b11111111;
		16'b1001010010111001: data <= 8'b11111111;
		16'b1001010010111010: data <= 8'b11111111;
		16'b1001010010111011: data <= 8'b11111111;
		16'b1001010010111100: data <= 8'b11111111;
		16'b1001010010111101: data <= 8'b11111111;
		16'b1001010010111110: data <= 8'b11111111;
		16'b1001010010111111: data <= 8'b11111111;
		16'b1001010011000000: data <= 8'b11111111;
		16'b1001010011000001: data <= 8'b11111111;
		16'b1001010011000010: data <= 8'b11111111;
		16'b1001010011000011: data <= 8'b11111111;
		16'b1001010011000100: data <= 8'b11111111;
		16'b1001010011000101: data <= 8'b11111111;
		16'b1001010011000110: data <= 8'b11111111;
		16'b1001010011000111: data <= 8'b11111111;
		16'b1001010011001000: data <= 8'b11111111;
		16'b1001010011001001: data <= 8'b11111111;
		16'b1001010011001010: data <= 8'b11111111;
		16'b1001010011001011: data <= 8'b11111111;
		16'b1001010011001100: data <= 8'b11111111;
		16'b1001010011001101: data <= 8'b11111111;
		16'b1001010011001110: data <= 8'b11111111;
		16'b1001010011001111: data <= 8'b11111111;
		16'b1001010011010000: data <= 8'b11111111;
		16'b1001010011010001: data <= 8'b11111111;
		16'b1001010011010010: data <= 8'b11111111;
		16'b1001010011010011: data <= 8'b11111111;
		16'b1001010011010100: data <= 8'b11111111;
		16'b1001010011010101: data <= 8'b11111111;
		16'b1001010011010110: data <= 8'b11111111;
		16'b1001010011010111: data <= 8'b11111111;
		16'b1001010011011000: data <= 8'b11111111;
		16'b1001010011011001: data <= 8'b11111111;
		16'b1001010011011010: data <= 8'b11111111;
		16'b1001010011011011: data <= 8'b11111111;
		16'b1001010011011100: data <= 8'b11111111;
		16'b1001010011011101: data <= 8'b11111111;
		16'b1001010011011110: data <= 8'b11111111;
		16'b1001010011011111: data <= 8'b11111111;
		16'b1001010011100000: data <= 8'b11111111;
		16'b1001010011100001: data <= 8'b11111111;
		16'b1001010011100010: data <= 8'b11111111;
		16'b1001010011100011: data <= 8'b11111111;
		16'b1001010011100100: data <= 8'b11111111;
		16'b1001010011100101: data <= 8'b11111111;
		16'b1001010011100110: data <= 8'b11111111;
		16'b1001010011100111: data <= 8'b11111111;
		16'b1001010011101000: data <= 8'b11111111;
		16'b1001010011101001: data <= 8'b11111111;
		16'b1001010011101010: data <= 8'b11111111;
		16'b1001010011101011: data <= 8'b11111111;
		16'b1001010011101100: data <= 8'b11111111;
		16'b1001010011101101: data <= 8'b11111111;
		16'b1001010011101110: data <= 8'b11111111;
		16'b1001010011101111: data <= 8'b11111111;
		16'b1001010011110000: data <= 8'b11111111;
		16'b1001010011110001: data <= 8'b11111111;
		16'b1001010011110010: data <= 8'b11111111;
		16'b1001010011110011: data <= 8'b11111111;
		16'b1001010011110100: data <= 8'b11111111;
		16'b1001010011110101: data <= 8'b11111111;
		16'b1001010011110110: data <= 8'b11111111;
		16'b1001010011110111: data <= 8'b11111111;
		16'b1001010011111000: data <= 8'b11111111;
		16'b1001010011111001: data <= 8'b11111111;
		16'b1001010011111010: data <= 8'b11111111;
		16'b1001010011111011: data <= 8'b11111111;
		16'b1001010011111100: data <= 8'b11111111;
		16'b1001010011111101: data <= 8'b11111111;
		16'b1001010011111110: data <= 8'b11111111;
		16'b1001010011111111: data <= 8'b11111111;
		16'b1001010100000000: data <= 8'b11111111;
		16'b1001010100000001: data <= 8'b11111111;
		16'b1001010100000010: data <= 8'b11111111;
		16'b1001010100000011: data <= 8'b11111111;
		16'b1001010100000100: data <= 8'b11111111;
		16'b1001010100000101: data <= 8'b11111111;
		16'b1001010100000110: data <= 8'b11111111;
		16'b1001010100000111: data <= 8'b11111111;
		16'b1001010100001000: data <= 8'b11111111;
		16'b1001010100001001: data <= 8'b11111111;
		16'b1001010100001010: data <= 8'b11111111;
		16'b1001010100001011: data <= 8'b11111111;
		16'b1001010100001100: data <= 8'b11111111;
		16'b1001010100001101: data <= 8'b11111111;
		16'b1001010100001110: data <= 8'b11111111;
		16'b1001010100001111: data <= 8'b11111111;
		16'b1001010100010000: data <= 8'b11111111;
		16'b1001010100010001: data <= 8'b11111111;
		16'b1001010100010010: data <= 8'b11111111;
		16'b1001010100010011: data <= 8'b11111111;
		16'b1001010100010100: data <= 8'b11111111;
		16'b1001010100010101: data <= 8'b11111111;
		16'b1001010100010110: data <= 8'b11111111;
		16'b1001010100010111: data <= 8'b11111111;
		16'b1001010100011000: data <= 8'b11111111;
		16'b1001010100011001: data <= 8'b11111111;
		16'b1001010100011010: data <= 8'b11111111;
		16'b1001010100011011: data <= 8'b11111111;
		16'b1001010100011100: data <= 8'b11111111;
		16'b1001010100011101: data <= 8'b11111111;
		16'b1001010100011110: data <= 8'b11111111;
		16'b1001010100011111: data <= 8'b11111111;
		16'b1001010100100000: data <= 8'b11111111;
		16'b1001010100100001: data <= 8'b11111111;
		16'b1001010100100010: data <= 8'b11111111;
		16'b1001010100100011: data <= 8'b11111111;
		16'b1001010100100100: data <= 8'b11111111;
		16'b1001010100100101: data <= 8'b11111111;
		16'b1001010100100110: data <= 8'b11111111;
		16'b1001010100100111: data <= 8'b11111111;
		16'b1001010100101000: data <= 8'b11111111;
		16'b1001010100101001: data <= 8'b11111111;
		16'b1001010100101010: data <= 8'b11111111;
		16'b1001010100101011: data <= 8'b11111111;
		16'b1001010100101100: data <= 8'b11111111;
		16'b1001010100101101: data <= 8'b11111111;
		16'b1001010100101110: data <= 8'b11111111;
		16'b1001010100101111: data <= 8'b11111111;
		16'b1001010100110000: data <= 8'b11111111;
		16'b1001010100110001: data <= 8'b11111111;
		16'b1001010100110010: data <= 8'b11111111;
		16'b1001010100110011: data <= 8'b11111111;
		16'b1001010100110100: data <= 8'b11111111;
		16'b1001010100110101: data <= 8'b11111111;
		16'b1001010100110110: data <= 8'b11111111;
		16'b1001010100110111: data <= 8'b11111111;
		16'b1001010100111000: data <= 8'b11111111;
		16'b1001010100111001: data <= 8'b11111111;
		16'b1001010100111010: data <= 8'b11111111;
		16'b1001010100111011: data <= 8'b11111111;
		16'b1001010100111100: data <= 8'b11111111;
		16'b1001010100111101: data <= 8'b11111111;
		16'b1001010100111110: data <= 8'b11111111;
		16'b1001010100111111: data <= 8'b11111111;
		16'b1001010101000000: data <= 8'b11111111;
		16'b1001010101000001: data <= 8'b11111111;
		16'b1001010101000010: data <= 8'b11111111;
		16'b1001010101000011: data <= 8'b11111111;
		16'b1001010101000100: data <= 8'b11111111;
		16'b1001010101000101: data <= 8'b11111111;
		16'b1001010101000110: data <= 8'b11111111;
		16'b1001010101000111: data <= 8'b11111111;
		16'b1001010101001000: data <= 8'b11111111;
		16'b1001010101001001: data <= 8'b11111111;
		16'b1001010101001010: data <= 8'b11111111;
		16'b1001010101001011: data <= 8'b11111111;
		16'b1001010101001100: data <= 8'b11111111;
		16'b1001010101001101: data <= 8'b11111111;
		16'b1001010101001110: data <= 8'b11111111;
		16'b1001010101001111: data <= 8'b11111111;
		16'b1001010101010000: data <= 8'b11111111;
		16'b1001010101010001: data <= 8'b11111111;
		16'b1001010101010010: data <= 8'b11111111;
		16'b1001010101010011: data <= 8'b11111111;
		16'b1001010101010100: data <= 8'b11111111;
		16'b1001010101010101: data <= 8'b11111111;
		16'b1001010101010110: data <= 8'b11111111;
		16'b1001010101010111: data <= 8'b11111111;
		16'b1001010101011000: data <= 8'b11111111;
		16'b1001010101011001: data <= 8'b11111111;
		16'b1001010101011010: data <= 8'b11111111;
		16'b1001010101011011: data <= 8'b11111111;
		16'b1001010101011100: data <= 8'b11111111;
		16'b1001010101011101: data <= 8'b11111111;
		16'b1001010101011110: data <= 8'b11111111;
		16'b1001010101011111: data <= 8'b11111111;
		16'b1001010101100000: data <= 8'b11111111;
		16'b1001010101100001: data <= 8'b11111111;
		16'b1001010101100010: data <= 8'b11111111;
		16'b1001010101100011: data <= 8'b11111111;
		16'b1001010101100100: data <= 8'b11111111;
		16'b1001010101100101: data <= 8'b11111111;
		16'b1001010101100110: data <= 8'b11111111;
		16'b1001010101100111: data <= 8'b11111111;
		16'b1001010101101000: data <= 8'b11111111;
		16'b1001010101101001: data <= 8'b11111111;
		16'b1001010101101010: data <= 8'b11111111;
		16'b1001010101101011: data <= 8'b11111111;
		16'b1001010101101100: data <= 8'b11111111;
		16'b1001010101101101: data <= 8'b11111111;
		16'b1001010101101110: data <= 8'b11111111;
		16'b1001010101101111: data <= 8'b11111111;
		16'b1001010101110000: data <= 8'b11111111;
		16'b1001010101110001: data <= 8'b11111111;
		16'b1001010101110010: data <= 8'b11111111;
		16'b1001010101110011: data <= 8'b11111111;
		16'b1001010101110100: data <= 8'b11111111;
		16'b1001010101110101: data <= 8'b11111111;
		16'b1001010101110110: data <= 8'b11111111;
		16'b1001010101110111: data <= 8'b11111111;
		16'b1001010101111000: data <= 8'b11111111;
		16'b1001010101111001: data <= 8'b11111111;
		16'b1001010101111010: data <= 8'b11111111;
		16'b1001010101111011: data <= 8'b11111111;
		16'b1001010101111100: data <= 8'b11111111;
		16'b1001010101111101: data <= 8'b11111111;
		16'b1001010101111110: data <= 8'b11111111;
		16'b1001010101111111: data <= 8'b11111111;
		16'b1001010110000000: data <= 8'b11111111;
		16'b1001010110000001: data <= 8'b11111111;
		16'b1001010110000010: data <= 8'b11111111;
		16'b1001010110000011: data <= 8'b11111111;
		16'b1001010110000100: data <= 8'b11111111;
		16'b1001010110000101: data <= 8'b11111111;
		16'b1001010110000110: data <= 8'b11111111;
		16'b1001010110000111: data <= 8'b11111111;
		16'b1001010110001000: data <= 8'b11111111;
		16'b1001010110001001: data <= 8'b11111111;
		16'b1001010110001010: data <= 8'b11111111;
		16'b1001010110001011: data <= 8'b11111111;
		16'b1001010110001100: data <= 8'b11111111;
		16'b1001010110001101: data <= 8'b11111111;
		16'b1001010110001110: data <= 8'b11111111;
		16'b1001010110001111: data <= 8'b11111111;
		16'b1001010110010000: data <= 8'b11111111;
		16'b1001010110010001: data <= 8'b11111111;
		16'b1001010110010010: data <= 8'b11111111;
		16'b1001010110010011: data <= 8'b11111111;
		16'b1001010110010100: data <= 8'b11111111;
		16'b1001010110010101: data <= 8'b11111111;
		16'b1001010110010110: data <= 8'b11111111;
		16'b1001010110010111: data <= 8'b11111111;
		16'b1001010110011000: data <= 8'b11111111;
		16'b1001010110011001: data <= 8'b11111111;
		16'b1001010110011010: data <= 8'b11111111;
		16'b1001010110011011: data <= 8'b11111111;
		16'b1001010110011100: data <= 8'b11111111;
		16'b1001010110011101: data <= 8'b11111111;
		16'b1001010110011110: data <= 8'b11111111;
		16'b1001010110011111: data <= 8'b11111111;
		16'b1001010110100000: data <= 8'b11111111;
		16'b1001010110100001: data <= 8'b11111111;
		16'b1001010110100010: data <= 8'b11111111;
		16'b1001010110100011: data <= 8'b11111111;
		16'b1001010110100100: data <= 8'b11111111;
		16'b1001010110100101: data <= 8'b11111111;
		16'b1001010110100110: data <= 8'b11111111;
		16'b1001010110100111: data <= 8'b11111111;
		16'b1001010110101000: data <= 8'b11111111;
		16'b1001010110101001: data <= 8'b11111111;
		16'b1001010110101010: data <= 8'b11111111;
		16'b1001010110101011: data <= 8'b11111111;
		16'b1001010110101100: data <= 8'b11111111;
		16'b1001010110101101: data <= 8'b11111111;
		16'b1001010110101110: data <= 8'b11111111;
		16'b1001010110101111: data <= 8'b11111111;
		16'b1001010110110000: data <= 8'b11111111;
		16'b1001010110110001: data <= 8'b11111111;
		16'b1001010110110010: data <= 8'b11111111;
		16'b1001010110110011: data <= 8'b11111111;
		16'b1001010110110100: data <= 8'b11111111;
		16'b1001010110110101: data <= 8'b11111111;
		16'b1001010110110110: data <= 8'b11111111;
		16'b1001010110110111: data <= 8'b11111111;
		16'b1001010110111000: data <= 8'b11111111;
		16'b1001010110111001: data <= 8'b11111111;
		16'b1001010110111010: data <= 8'b11111111;
		16'b1001010110111011: data <= 8'b11111111;
		16'b1001010110111100: data <= 8'b11111111;
		16'b1001010110111101: data <= 8'b11111111;
		16'b1001010110111110: data <= 8'b11111111;
		16'b1001010110111111: data <= 8'b11111111;
		16'b1001010111000000: data <= 8'b11111111;
		16'b1001010111000001: data <= 8'b11111111;
		16'b1001010111000010: data <= 8'b11111111;
		16'b1001010111000011: data <= 8'b11111111;
		16'b1001010111000100: data <= 8'b11111111;
		16'b1001010111000101: data <= 8'b11111111;
		16'b1001010111000110: data <= 8'b11111111;
		16'b1001010111000111: data <= 8'b11111111;
		16'b1001010111001000: data <= 8'b11111111;
		16'b1001010111001001: data <= 8'b11111111;
		16'b1001010111001010: data <= 8'b11111111;
		16'b1001010111001011: data <= 8'b11111111;
		16'b1001010111001100: data <= 8'b11111111;
		16'b1001010111001101: data <= 8'b11111111;
		16'b1001010111001110: data <= 8'b11111111;
		16'b1001010111001111: data <= 8'b11111111;
		16'b1001010111010000: data <= 8'b11111111;
		16'b1001010111010001: data <= 8'b11111111;
		16'b1001010111010010: data <= 8'b11111111;
		16'b1001010111010011: data <= 8'b11111111;
		16'b1001010111010100: data <= 8'b11111111;
		16'b1001010111010101: data <= 8'b11111111;
		16'b1001010111010110: data <= 8'b11111111;
		16'b1001010111010111: data <= 8'b11111111;
		16'b1001010111011000: data <= 8'b11111111;
		16'b1001010111011001: data <= 8'b11111111;
		16'b1001010111011010: data <= 8'b11111111;
		16'b1001010111011011: data <= 8'b11111111;
		16'b1001010111011100: data <= 8'b11111111;
		16'b1001010111011101: data <= 8'b11111111;
		16'b1001010111011110: data <= 8'b11111111;
		16'b1001010111011111: data <= 8'b11111111;
		16'b1001010111100000: data <= 8'b11111111;
		16'b1001010111100001: data <= 8'b11111111;
		16'b1001010111100010: data <= 8'b11111111;
		16'b1001010111100011: data <= 8'b11111111;
		16'b1001010111100100: data <= 8'b11111111;
		16'b1001010111100101: data <= 8'b11111111;
		16'b1001010111100110: data <= 8'b11111111;
		16'b1001010111100111: data <= 8'b11111111;
		16'b1001010111101000: data <= 8'b11111111;
		16'b1001010111101001: data <= 8'b11111111;
		16'b1001010111101010: data <= 8'b11111111;
		16'b1001010111101011: data <= 8'b11111111;
		16'b1001010111101100: data <= 8'b11111111;
		16'b1001010111101101: data <= 8'b11111111;
		16'b1001010111101110: data <= 8'b11111111;
		16'b1001010111101111: data <= 8'b11111111;
		16'b1001010111110000: data <= 8'b11111111;
		16'b1001010111110001: data <= 8'b11111111;
		16'b1001010111110010: data <= 8'b11111111;
		16'b1001010111110011: data <= 8'b11111111;
		16'b1001010111110100: data <= 8'b11111111;
		16'b1001010111110101: data <= 8'b11111111;
		16'b1001010111110110: data <= 8'b11111111;
		16'b1001010111110111: data <= 8'b11111111;
		16'b1001010111111000: data <= 8'b11111111;
		16'b1001010111111001: data <= 8'b11111111;
		16'b1001010111111010: data <= 8'b11111111;
		16'b1001010111111011: data <= 8'b11111111;
		16'b1001010111111100: data <= 8'b11111111;
		16'b1001010111111101: data <= 8'b11111111;
		16'b1001010111111110: data <= 8'b11111111;
		16'b1001010111111111: data <= 8'b11111111;
		16'b1001011000000000: data <= 8'b11111111;
		16'b1001011000000001: data <= 8'b11111111;
		16'b1001011000000010: data <= 8'b11111111;
		16'b1001011000000011: data <= 8'b11111111;
		16'b1001011000000100: data <= 8'b11111111;
		16'b1001011000000101: data <= 8'b11111111;
		16'b1001011000000110: data <= 8'b11111111;
		16'b1001011000000111: data <= 8'b11111111;
		16'b1001011000001000: data <= 8'b11111111;
		16'b1001011000001001: data <= 8'b11111111;
		16'b1001011000001010: data <= 8'b11111111;
		16'b1001011000001011: data <= 8'b11111111;
		16'b1001011000001100: data <= 8'b11111111;
		16'b1001011000001101: data <= 8'b11111111;
		16'b1001011000001110: data <= 8'b11111111;
		16'b1001011000001111: data <= 8'b11111111;
		16'b1001011000010000: data <= 8'b11111111;
		16'b1001011000010001: data <= 8'b11111111;
		16'b1001011000010010: data <= 8'b11111111;
		16'b1001011000010011: data <= 8'b11111111;
		16'b1001011000010100: data <= 8'b11111111;
		16'b1001011000010101: data <= 8'b11111111;
		16'b1001011000010110: data <= 8'b11111111;
		16'b1001011000010111: data <= 8'b11111111;
		16'b1001011000011000: data <= 8'b11111111;
		16'b1001011000011001: data <= 8'b11111111;
		16'b1001011000011010: data <= 8'b11111111;
		16'b1001011000011011: data <= 8'b11111111;
		16'b1001011000011100: data <= 8'b11111111;
		16'b1001011000011101: data <= 8'b11111111;
		16'b1001011000011110: data <= 8'b11111111;
		16'b1001011000011111: data <= 8'b11111111;
		16'b1001011000100000: data <= 8'b11111111;
		16'b1001011000100001: data <= 8'b11111111;
		16'b1001011000100010: data <= 8'b11111111;
		16'b1001011000100011: data <= 8'b11111111;
		16'b1001011000100100: data <= 8'b11111111;
		16'b1001011000100101: data <= 8'b11111111;
		16'b1001011000100110: data <= 8'b11111111;
		16'b1001011000100111: data <= 8'b11111111;
		16'b1001011000101000: data <= 8'b11111111;
		16'b1001011000101001: data <= 8'b11111111;
		16'b1001011000101010: data <= 8'b11111111;
		16'b1001011000101011: data <= 8'b11111111;
		16'b1001011000101100: data <= 8'b11111111;
		16'b1001011000101101: data <= 8'b11111111;
		16'b1001011000101110: data <= 8'b11111111;
		16'b1001011000101111: data <= 8'b11111111;
		16'b1001011000110000: data <= 8'b11111111;
		16'b1001011000110001: data <= 8'b11111111;
		16'b1001011000110010: data <= 8'b11111111;
		16'b1001011000110011: data <= 8'b11111111;
		16'b1001011000110100: data <= 8'b11111111;
		16'b1001011000110101: data <= 8'b11111111;
		16'b1001011000110110: data <= 8'b11111111;
		16'b1001011000110111: data <= 8'b11111111;
		16'b1001011000111000: data <= 8'b11111111;
		16'b1001011000111001: data <= 8'b11111111;
		16'b1001011000111010: data <= 8'b11111111;
		16'b1001011000111011: data <= 8'b11111111;
		16'b1001011000111100: data <= 8'b11111111;
		16'b1001011000111101: data <= 8'b11111111;
		16'b1001011000111110: data <= 8'b11111111;
		16'b1001011000111111: data <= 8'b11111111;
		16'b1001011001000000: data <= 8'b11111111;
		16'b1001011001000001: data <= 8'b11111111;
		16'b1001011001000010: data <= 8'b11111111;
		16'b1001011001000011: data <= 8'b11111111;
		16'b1001011001000100: data <= 8'b11111111;
		16'b1001011001000101: data <= 8'b11111111;
		16'b1001011001000110: data <= 8'b11111111;
		16'b1001011001000111: data <= 8'b11111111;
		16'b1001011001001000: data <= 8'b11111111;
		16'b1001011001001001: data <= 8'b11111111;
		16'b1001011001001010: data <= 8'b11111111;
		16'b1001011001001011: data <= 8'b11111111;
		16'b1001011001001100: data <= 8'b11111111;
		16'b1001011001001101: data <= 8'b11111111;
		16'b1001011001001110: data <= 8'b11111111;
		16'b1001011001001111: data <= 8'b11111111;
		16'b1001011001010000: data <= 8'b11111111;
		16'b1001011001010001: data <= 8'b11111111;
		16'b1001011001010010: data <= 8'b11111111;
		16'b1001011001010011: data <= 8'b11111111;
		16'b1001011001010100: data <= 8'b11111111;
		16'b1001011001010101: data <= 8'b11111111;
		16'b1001011001010110: data <= 8'b11111111;
		16'b1001011001010111: data <= 8'b11111111;
		16'b1001011001011000: data <= 8'b11111111;
		16'b1001011001011001: data <= 8'b11111111;
		16'b1001011001011010: data <= 8'b11111111;
		16'b1001011001011011: data <= 8'b11111111;
		16'b1001011001011100: data <= 8'b11111111;
		16'b1001011001011101: data <= 8'b11111111;
		16'b1001011001011110: data <= 8'b11111111;
		16'b1001011001011111: data <= 8'b11111111;
		16'b1001011001100000: data <= 8'b11111111;
		16'b1001011001100001: data <= 8'b11111111;
		16'b1001011001100010: data <= 8'b11111111;
		16'b1001011001100011: data <= 8'b11111111;
		16'b1001011001100100: data <= 8'b11111111;
		16'b1001011001100101: data <= 8'b11111111;
		16'b1001011001100110: data <= 8'b11111111;
		16'b1001011001100111: data <= 8'b11111111;
		16'b1001011001101000: data <= 8'b11111111;
		16'b1001011001101001: data <= 8'b11111111;
		16'b1001011001101010: data <= 8'b11111111;
		16'b1001011001101011: data <= 8'b11111111;
		16'b1001011001101100: data <= 8'b11111111;
		16'b1001011001101101: data <= 8'b11111111;
		16'b1001011001101110: data <= 8'b11111111;
		16'b1001011001101111: data <= 8'b11111111;
		16'b1001011001110000: data <= 8'b11111111;
		16'b1001011001110001: data <= 8'b11111111;
		16'b1001011001110010: data <= 8'b11111111;
		16'b1001011001110011: data <= 8'b11111111;
		16'b1001011001110100: data <= 8'b11111111;
		16'b1001011001110101: data <= 8'b11111111;
		16'b1001011001110110: data <= 8'b11111111;
		16'b1001011001110111: data <= 8'b11111111;
		16'b1001011001111000: data <= 8'b11111111;
		16'b1001011001111001: data <= 8'b11111111;
		16'b1001011001111010: data <= 8'b11111111;
		16'b1001011001111011: data <= 8'b11111111;
		16'b1001011001111100: data <= 8'b11111111;
		16'b1001011001111101: data <= 8'b11111111;
		16'b1001011001111110: data <= 8'b11111111;
		16'b1001011001111111: data <= 8'b11111111;
		16'b1001011010000000: data <= 8'b11111111;
		16'b1001011010000001: data <= 8'b11111111;
		16'b1001011010000010: data <= 8'b11111111;
		16'b1001011010000011: data <= 8'b11111111;
		16'b1001011010000100: data <= 8'b11111111;
		16'b1001011010000101: data <= 8'b11111111;
		16'b1001011010000110: data <= 8'b11111111;
		16'b1001011010000111: data <= 8'b11111111;
		16'b1001011010001000: data <= 8'b11111111;
		16'b1001011010001001: data <= 8'b11111111;
		16'b1001011010001010: data <= 8'b11111111;
		16'b1001011010001011: data <= 8'b11111111;
		16'b1001011010001100: data <= 8'b11111111;
		16'b1001011010001101: data <= 8'b11111111;
		16'b1001011010001110: data <= 8'b11111111;
		16'b1001011010001111: data <= 8'b11111111;
		16'b1001011010010000: data <= 8'b11111111;
		16'b1001011010010001: data <= 8'b11111111;
		16'b1001011010010010: data <= 8'b11111111;
		16'b1001011010010011: data <= 8'b11111111;
		16'b1001011010010100: data <= 8'b11111111;
		16'b1001011010010101: data <= 8'b11111111;
		16'b1001011010010110: data <= 8'b11111111;
		16'b1001011010010111: data <= 8'b11111111;
		16'b1001011010011000: data <= 8'b11111111;
		16'b1001011010011001: data <= 8'b11111111;
		16'b1001011010011010: data <= 8'b11111111;
		16'b1001011010011011: data <= 8'b11111111;
		16'b1001011010011100: data <= 8'b11111111;
		16'b1001011010011101: data <= 8'b11111111;
		16'b1001011010011110: data <= 8'b11111111;
		16'b1001011010011111: data <= 8'b11111111;
		16'b1001011010100000: data <= 8'b11111111;
		16'b1001011010100001: data <= 8'b11111111;
		16'b1001011010100010: data <= 8'b11111111;
		16'b1001011010100011: data <= 8'b11111111;
		16'b1001011010100100: data <= 8'b11111111;
		16'b1001011010100101: data <= 8'b11111111;
		16'b1001011010100110: data <= 8'b11111111;
		16'b1001011010100111: data <= 8'b11111111;
		16'b1001011010101000: data <= 8'b11111111;
		16'b1001011010101001: data <= 8'b11111111;
		16'b1001011010101010: data <= 8'b11111111;
		16'b1001011010101011: data <= 8'b11111111;
		16'b1001011010101100: data <= 8'b11111111;
		16'b1001011010101101: data <= 8'b11111111;
		16'b1001011010101110: data <= 8'b11111111;
		16'b1001011010101111: data <= 8'b11111111;
		16'b1001011010110000: data <= 8'b11111111;
		16'b1001011010110001: data <= 8'b11111111;
		16'b1001011010110010: data <= 8'b11111111;
		16'b1001011010110011: data <= 8'b11111111;
		16'b1001011010110100: data <= 8'b11111111;
		16'b1001011010110101: data <= 8'b11111111;
		16'b1001011010110110: data <= 8'b11111111;
		16'b1001011010110111: data <= 8'b11111111;
		16'b1001011010111000: data <= 8'b11111111;
		16'b1001011010111001: data <= 8'b11111111;
		16'b1001011010111010: data <= 8'b11111111;
		16'b1001011010111011: data <= 8'b11111111;
		16'b1001011010111100: data <= 8'b11111111;
		16'b1001011010111101: data <= 8'b11111111;
		16'b1001011010111110: data <= 8'b11111111;
		16'b1001011010111111: data <= 8'b11111111;
		16'b1001011011000000: data <= 8'b11111111;
		16'b1001011011000001: data <= 8'b11111111;
		16'b1001011011000010: data <= 8'b11111111;
		16'b1001011011000011: data <= 8'b11111111;
		16'b1001011011000100: data <= 8'b11111111;
		16'b1001011011000101: data <= 8'b11111111;
		16'b1001011011000110: data <= 8'b11111111;
		16'b1001011011000111: data <= 8'b11111111;
		16'b1001011011001000: data <= 8'b11111111;
		16'b1001011011001001: data <= 8'b11111111;
		16'b1001011011001010: data <= 8'b11111111;
		16'b1001011011001011: data <= 8'b11111111;
		16'b1001011011001100: data <= 8'b11111111;
		16'b1001011011001101: data <= 8'b11111111;
		16'b1001011011001110: data <= 8'b11111111;
		16'b1001011011001111: data <= 8'b11111111;
		16'b1001011011010000: data <= 8'b11111111;
		16'b1001011011010001: data <= 8'b11111111;
		16'b1001011011010010: data <= 8'b11111111;
		16'b1001011011010011: data <= 8'b11111111;
		16'b1001011011010100: data <= 8'b11111111;
		16'b1001011011010101: data <= 8'b11111111;
		16'b1001011011010110: data <= 8'b11111111;
		16'b1001011011010111: data <= 8'b11111111;
		16'b1001011011011000: data <= 8'b11111111;
		16'b1001011011011001: data <= 8'b11111111;
		16'b1001011011011010: data <= 8'b11111111;
		16'b1001011011011011: data <= 8'b11111111;
		16'b1001011011011100: data <= 8'b11111111;
		16'b1001011011011101: data <= 8'b11111111;
		16'b1001011011011110: data <= 8'b11111111;
		16'b1001011011011111: data <= 8'b11111111;
		16'b1001011011100000: data <= 8'b11111111;
		16'b1001011011100001: data <= 8'b11111111;
		16'b1001011011100010: data <= 8'b11111111;
		16'b1001011011100011: data <= 8'b11111111;
		16'b1001011011100100: data <= 8'b11111111;
		16'b1001011011100101: data <= 8'b11111111;
		16'b1001011011100110: data <= 8'b11111111;
		16'b1001011011100111: data <= 8'b11111111;
		16'b1001011011101000: data <= 8'b11111111;
		16'b1001011011101001: data <= 8'b11111111;
		16'b1001011011101010: data <= 8'b11111111;
		16'b1001011011101011: data <= 8'b11111111;
		16'b1001011011101100: data <= 8'b11111111;
		16'b1001011011101101: data <= 8'b11111111;
		16'b1001011011101110: data <= 8'b11111111;
		16'b1001011011101111: data <= 8'b11111111;
		16'b1001011011110000: data <= 8'b11111111;
		16'b1001011011110001: data <= 8'b11111111;
		16'b1001011011110010: data <= 8'b11111111;
		16'b1001011011110011: data <= 8'b11111111;
		16'b1001011011110100: data <= 8'b11111111;
		16'b1001011011110101: data <= 8'b11111111;
		16'b1001011011110110: data <= 8'b11111111;
		16'b1001011011110111: data <= 8'b11111111;
		16'b1001011011111000: data <= 8'b11111111;
		16'b1001011011111001: data <= 8'b11111111;
		16'b1001011011111010: data <= 8'b11111111;
		16'b1001011011111011: data <= 8'b11111111;
		16'b1001011011111100: data <= 8'b11111111;
		16'b1001011011111101: data <= 8'b11111111;
		16'b1001011011111110: data <= 8'b11111111;
		16'b1001011011111111: data <= 8'b11111111;
		16'b1001011100000000: data <= 8'b11111111;
		16'b1001011100000001: data <= 8'b11111111;
		16'b1001011100000010: data <= 8'b11111111;
		16'b1001011100000011: data <= 8'b11111111;
		16'b1001011100000100: data <= 8'b11111111;
		16'b1001011100000101: data <= 8'b11111111;
		16'b1001011100000110: data <= 8'b11111111;
		16'b1001011100000111: data <= 8'b11111111;
		16'b1001011100001000: data <= 8'b11111111;
		16'b1001011100001001: data <= 8'b11111111;
		16'b1001011100001010: data <= 8'b11111111;
		16'b1001011100001011: data <= 8'b11111111;
		16'b1001011100001100: data <= 8'b11111111;
		16'b1001011100001101: data <= 8'b11111111;
		16'b1001011100001110: data <= 8'b11111111;
		16'b1001011100001111: data <= 8'b11111111;
		16'b1001011100010000: data <= 8'b11111111;
		16'b1001011100010001: data <= 8'b11111111;
		16'b1001011100010010: data <= 8'b11111111;
		16'b1001011100010011: data <= 8'b11111111;
		16'b1001011100010100: data <= 8'b11111111;
		16'b1001011100010101: data <= 8'b11111111;
		16'b1001011100010110: data <= 8'b11111111;
		16'b1001011100010111: data <= 8'b11111111;
		16'b1001011100011000: data <= 8'b11111111;
		16'b1001011100011001: data <= 8'b11111111;
		16'b1001011100011010: data <= 8'b11111111;
		16'b1001011100011011: data <= 8'b11111111;
		16'b1001011100011100: data <= 8'b11111111;
		16'b1001011100011101: data <= 8'b11111111;
		16'b1001011100011110: data <= 8'b11111111;
		16'b1001011100011111: data <= 8'b11111111;
		16'b1001011100100000: data <= 8'b11111111;
		16'b1001011100100001: data <= 8'b11111111;
		16'b1001011100100010: data <= 8'b11111111;
		16'b1001011100100011: data <= 8'b11111111;
		16'b1001011100100100: data <= 8'b11111111;
		16'b1001011100100101: data <= 8'b11111111;
		16'b1001011100100110: data <= 8'b11111111;
		16'b1001011100100111: data <= 8'b11111111;
		16'b1001011100101000: data <= 8'b11111111;
		16'b1001011100101001: data <= 8'b11111111;
		16'b1001011100101010: data <= 8'b11111111;
		16'b1001011100101011: data <= 8'b11111111;
		16'b1001011100101100: data <= 8'b11111111;
		16'b1001011100101101: data <= 8'b11111111;
		16'b1001011100101110: data <= 8'b11111111;
		16'b1001011100101111: data <= 8'b11111111;
		16'b1001011100110000: data <= 8'b11111111;
		16'b1001011100110001: data <= 8'b11111111;
		16'b1001011100110010: data <= 8'b11111111;
		16'b1001011100110011: data <= 8'b11111111;
		16'b1001011100110100: data <= 8'b11111111;
		16'b1001011100110101: data <= 8'b11111111;
		16'b1001011100110110: data <= 8'b11111111;
		16'b1001011100110111: data <= 8'b11111111;
		16'b1001011100111000: data <= 8'b11111111;
		16'b1001011100111001: data <= 8'b11111111;
		16'b1001011100111010: data <= 8'b11111111;
		16'b1001011100111011: data <= 8'b11111111;
		16'b1001011100111100: data <= 8'b11111111;
		16'b1001011100111101: data <= 8'b11111111;
		16'b1001011100111110: data <= 8'b11111111;
		16'b1001011100111111: data <= 8'b11111111;
		16'b1001011101000000: data <= 8'b11111111;
		16'b1001011101000001: data <= 8'b11111111;
		16'b1001011101000010: data <= 8'b11111111;
		16'b1001011101000011: data <= 8'b11111111;
		16'b1001011101000100: data <= 8'b11111111;
		16'b1001011101000101: data <= 8'b11111111;
		16'b1001011101000110: data <= 8'b11111111;
		16'b1001011101000111: data <= 8'b11111111;
		16'b1001011101001000: data <= 8'b11111111;
		16'b1001011101001001: data <= 8'b11111111;
		16'b1001011101001010: data <= 8'b11111111;
		16'b1001011101001011: data <= 8'b11111111;
		16'b1001011101001100: data <= 8'b11111111;
		16'b1001011101001101: data <= 8'b11111111;
		16'b1001011101001110: data <= 8'b11111111;
		16'b1001011101001111: data <= 8'b11111111;
		16'b1001011101010000: data <= 8'b11111111;
		16'b1001011101010001: data <= 8'b11111111;
		16'b1001011101010010: data <= 8'b11111111;
		16'b1001011101010011: data <= 8'b11111111;
		16'b1001011101010100: data <= 8'b11111111;
		16'b1001011101010101: data <= 8'b11111111;
		16'b1001011101010110: data <= 8'b11111111;
		16'b1001011101010111: data <= 8'b11111111;
		16'b1001011101011000: data <= 8'b11111111;
		16'b1001011101011001: data <= 8'b11111111;
		16'b1001011101011010: data <= 8'b11111111;
		16'b1001011101011011: data <= 8'b11111111;
		16'b1001011101011100: data <= 8'b11111111;
		16'b1001011101011101: data <= 8'b11111111;
		16'b1001011101011110: data <= 8'b11111111;
		16'b1001011101011111: data <= 8'b11111111;
		16'b1001011101100000: data <= 8'b11111111;
		16'b1001011101100001: data <= 8'b11111111;
		16'b1001011101100010: data <= 8'b11111111;
		16'b1001011101100011: data <= 8'b11111111;
		16'b1001011101100100: data <= 8'b11111111;
		16'b1001011101100101: data <= 8'b11111111;
		16'b1001011101100110: data <= 8'b11111111;
		16'b1001011101100111: data <= 8'b11111111;
		16'b1001011101101000: data <= 8'b11111111;
		16'b1001011101101001: data <= 8'b11111111;
		16'b1001011101101010: data <= 8'b11111111;
		16'b1001011101101011: data <= 8'b11111111;
		16'b1001011101101100: data <= 8'b11111111;
		16'b1001011101101101: data <= 8'b11111111;
		16'b1001011101101110: data <= 8'b11111111;
		16'b1001011101101111: data <= 8'b11111111;
		16'b1001011101110000: data <= 8'b11111111;
		16'b1001011101110001: data <= 8'b11111111;
		16'b1001011101110010: data <= 8'b11111111;
		16'b1001011101110011: data <= 8'b11111111;
		16'b1001011101110100: data <= 8'b11111111;
		16'b1001011101110101: data <= 8'b11111111;
		16'b1001011101110110: data <= 8'b11111111;
		16'b1001011101110111: data <= 8'b11111111;
		16'b1001011101111000: data <= 8'b11111111;
		16'b1001011101111001: data <= 8'b11111111;
		16'b1001011101111010: data <= 8'b11111111;
		16'b1001011101111011: data <= 8'b11111111;
		16'b1001011101111100: data <= 8'b11111111;
		16'b1001011101111101: data <= 8'b11111111;
		16'b1001011101111110: data <= 8'b11111111;
		16'b1001011101111111: data <= 8'b11111111;
		16'b1001011110000000: data <= 8'b11111111;
		16'b1001011110000001: data <= 8'b11111111;
		16'b1001011110000010: data <= 8'b11111111;
		16'b1001011110000011: data <= 8'b11111111;
		16'b1001011110000100: data <= 8'b11111111;
		16'b1001011110000101: data <= 8'b11111111;
		16'b1001011110000110: data <= 8'b11111111;
		16'b1001011110000111: data <= 8'b11111111;
		16'b1001011110001000: data <= 8'b11111111;
		16'b1001011110001001: data <= 8'b11111111;
		16'b1001011110001010: data <= 8'b11111111;
		16'b1001011110001011: data <= 8'b11111111;
		16'b1001011110001100: data <= 8'b11111111;
		16'b1001011110001101: data <= 8'b11111111;
		16'b1001011110001110: data <= 8'b11111111;
		16'b1001011110001111: data <= 8'b11111111;
		16'b1001011110010000: data <= 8'b11111111;
		16'b1001011110010001: data <= 8'b11111111;
		16'b1001011110010010: data <= 8'b11111111;
		16'b1001011110010011: data <= 8'b11111111;
		16'b1001011110010100: data <= 8'b11111111;
		16'b1001011110010101: data <= 8'b11111111;
		16'b1001011110010110: data <= 8'b11111111;
		16'b1001011110010111: data <= 8'b11111111;
		16'b1001011110011000: data <= 8'b11111111;
		16'b1001011110011001: data <= 8'b11111111;
		16'b1001011110011010: data <= 8'b11111111;
		16'b1001011110011011: data <= 8'b11111111;
		16'b1001011110011100: data <= 8'b11111111;
		16'b1001011110011101: data <= 8'b11111111;
		16'b1001011110011110: data <= 8'b11111111;
		16'b1001011110011111: data <= 8'b11111111;
		16'b1001011110100000: data <= 8'b11111111;
		16'b1001011110100001: data <= 8'b11111111;
		16'b1001011110100010: data <= 8'b11111111;
		16'b1001011110100011: data <= 8'b11111111;
		16'b1001011110100100: data <= 8'b11111111;
		16'b1001011110100101: data <= 8'b11111111;
		16'b1001011110100110: data <= 8'b11111111;
		16'b1001011110100111: data <= 8'b11111111;
		16'b1001011110101000: data <= 8'b11111111;
		16'b1001011110101001: data <= 8'b11111111;
		16'b1001011110101010: data <= 8'b11111111;
		16'b1001011110101011: data <= 8'b11111111;
		16'b1001011110101100: data <= 8'b11111111;
		16'b1001011110101101: data <= 8'b11111111;
		16'b1001011110101110: data <= 8'b11111111;
		16'b1001011110101111: data <= 8'b11111111;
		16'b1001011110110000: data <= 8'b11111111;
		16'b1001011110110001: data <= 8'b11111111;
		16'b1001011110110010: data <= 8'b11111111;
		16'b1001011110110011: data <= 8'b11111111;
		16'b1001011110110100: data <= 8'b11111111;
		16'b1001011110110101: data <= 8'b11111111;
		16'b1001011110110110: data <= 8'b11111111;
		16'b1001011110110111: data <= 8'b11111111;
		16'b1001011110111000: data <= 8'b11111111;
		16'b1001011110111001: data <= 8'b11111111;
		16'b1001011110111010: data <= 8'b11111111;
		16'b1001011110111011: data <= 8'b11111111;
		16'b1001011110111100: data <= 8'b11111111;
		16'b1001011110111101: data <= 8'b11111111;
		16'b1001011110111110: data <= 8'b11111111;
		16'b1001011110111111: data <= 8'b11111111;
		16'b1001011111000000: data <= 8'b11111111;
		16'b1001011111000001: data <= 8'b11111111;
		16'b1001011111000010: data <= 8'b11111111;
		16'b1001011111000011: data <= 8'b11111111;
		16'b1001011111000100: data <= 8'b11111111;
		16'b1001011111000101: data <= 8'b11111111;
		16'b1001011111000110: data <= 8'b11111111;
		16'b1001011111000111: data <= 8'b11111111;
		16'b1001011111001000: data <= 8'b11111111;
		16'b1001011111001001: data <= 8'b11111111;
		16'b1001011111001010: data <= 8'b11111111;
		16'b1001011111001011: data <= 8'b11111111;
		16'b1001011111001100: data <= 8'b11111111;
		16'b1001011111001101: data <= 8'b11111111;
		16'b1001011111001110: data <= 8'b11111111;
		16'b1001011111001111: data <= 8'b11111111;
		16'b1001011111010000: data <= 8'b11111111;
		16'b1001011111010001: data <= 8'b11111111;
		16'b1001011111010010: data <= 8'b11111111;
		16'b1001011111010011: data <= 8'b11111111;
		16'b1001011111010100: data <= 8'b11111111;
		16'b1001011111010101: data <= 8'b11111111;
		16'b1001011111010110: data <= 8'b11111111;
		16'b1001011111010111: data <= 8'b11111111;
		16'b1001011111011000: data <= 8'b11111111;
		16'b1001011111011001: data <= 8'b11111111;
		16'b1001011111011010: data <= 8'b11111111;
		16'b1001011111011011: data <= 8'b11111111;
		16'b1001011111011100: data <= 8'b11111111;
		16'b1001011111011101: data <= 8'b11111111;
		16'b1001011111011110: data <= 8'b11111111;
		16'b1001011111011111: data <= 8'b11111111;
		16'b1001100000101110: data <= 8'b11111111;
		16'b1001100000101111: data <= 8'b11111111;
		16'b1001100000110000: data <= 8'b11111111;
		16'b1001100000110001: data <= 8'b11111111;
		16'b1001100001111110: data <= 8'b11111111;
		16'b1001100001111111: data <= 8'b11111111;
		16'b1001100010000000: data <= 8'b11111111;
		16'b1001100010000001: data <= 8'b11111111;
		16'b1001100100011110: data <= 8'b11111111;
		16'b1001100100011111: data <= 8'b11111111;
		16'b1001100100100000: data <= 8'b11111111;
		16'b1001100100100001: data <= 8'b11111111;
		16'b1001100101101110: data <= 8'b11111111;
		16'b1001100101101111: data <= 8'b11111111;
		16'b1001100101110000: data <= 8'b11111111;
		16'b1001100101110001: data <= 8'b11111111;
		16'b1001101000001110: data <= 8'b11111111;
		16'b1001101000001111: data <= 8'b11111111;
		16'b1001101000010000: data <= 8'b11111111;
		16'b1001101000010001: data <= 8'b11111111;
		16'b1001101001011110: data <= 8'b11111111;
		16'b1001101001011111: data <= 8'b11111111;
		16'b1001101001100000: data <= 8'b11111111;
		16'b1001101001100001: data <= 8'b11111111;
		16'b1001101011111110: data <= 8'b11111111;
		16'b1001101011111111: data <= 8'b11111111;
		16'b1001101100000000: data <= 8'b11111111;
		16'b1001101100000001: data <= 8'b11111111;
		16'b1001101101001110: data <= 8'b11111111;
		16'b1001101101001111: data <= 8'b11111111;
		16'b1001101101010000: data <= 8'b11111111;
		16'b1001101101010001: data <= 8'b11111111;
		16'b1001101111101110: data <= 8'b11111111;
		16'b1001101111101111: data <= 8'b11111111;
		16'b1001101111110000: data <= 8'b11111111;
		16'b1001101111110001: data <= 8'b11111111;
		16'b1001110000111110: data <= 8'b11111111;
		16'b1001110000111111: data <= 8'b11111111;
		16'b1001110001000000: data <= 8'b11111111;
		16'b1001110001000001: data <= 8'b11111111;
		16'b1001110011011110: data <= 8'b11111111;
		16'b1001110011011111: data <= 8'b11111111;
		16'b1001110011100000: data <= 8'b11111111;
		16'b1001110011100001: data <= 8'b11111111;
		16'b1001110100101110: data <= 8'b11111111;
		16'b1001110100101111: data <= 8'b11111111;
		16'b1001110100110000: data <= 8'b11111111;
		16'b1001110100110001: data <= 8'b11111111;
		16'b1001110111001110: data <= 8'b11111111;
		16'b1001110111001111: data <= 8'b11111111;
		16'b1001110111010000: data <= 8'b11111111;
		16'b1001110111010001: data <= 8'b11111111;
		16'b1001111000011110: data <= 8'b11111111;
		16'b1001111000011111: data <= 8'b11111111;
		16'b1001111000100000: data <= 8'b11111111;
		16'b1001111000100001: data <= 8'b11111111;
		16'b1001111010111110: data <= 8'b11111111;
		16'b1001111010111111: data <= 8'b11111111;
		16'b1001111011000000: data <= 8'b11111111;
		16'b1001111011000001: data <= 8'b11111111;
		16'b1001111100001110: data <= 8'b11111111;
		16'b1001111100001111: data <= 8'b11111111;
		16'b1001111100010000: data <= 8'b11111111;
		16'b1001111100010001: data <= 8'b11111111;
		16'b1001111110101110: data <= 8'b11111111;
		16'b1001111110101111: data <= 8'b11111111;
		16'b1001111110110000: data <= 8'b11111111;
		16'b1001111110110001: data <= 8'b11111111;
		16'b1001111111111110: data <= 8'b11111111;
		16'b1001111111111111: data <= 8'b11111111;
		16'b1010000000000000: data <= 8'b11111111;
		16'b1010000000000001: data <= 8'b11111111;
		16'b1010000010011110: data <= 8'b11111111;
		16'b1010000010011111: data <= 8'b11111111;
		16'b1010000010100000: data <= 8'b11111111;
		16'b1010000010100001: data <= 8'b11111111;
		16'b1010000011101110: data <= 8'b11111111;
		16'b1010000011101111: data <= 8'b11111111;
		16'b1010000011110000: data <= 8'b11111111;
		16'b1010000011110001: data <= 8'b11111111;
		16'b1010000110001110: data <= 8'b11111111;
		16'b1010000110001111: data <= 8'b11111111;
		16'b1010000110010000: data <= 8'b11111111;
		16'b1010000110010001: data <= 8'b11111111;
		16'b1010000111011110: data <= 8'b11111111;
		16'b1010000111011111: data <= 8'b11111111;
		16'b1010000111100000: data <= 8'b11111111;
		16'b1010000111100001: data <= 8'b11111111;
		16'b1010001001111110: data <= 8'b11111111;
		16'b1010001001111111: data <= 8'b11111111;
		16'b1010001010000000: data <= 8'b11111111;
		16'b1010001010000001: data <= 8'b11111111;
		16'b1010001011001110: data <= 8'b11111111;
		16'b1010001011001111: data <= 8'b11111111;
		16'b1010001011010000: data <= 8'b11111111;
		16'b1010001011010001: data <= 8'b11111111;
		16'b1010001101101110: data <= 8'b11111111;
		16'b1010001101101111: data <= 8'b11111111;
		16'b1010001101110000: data <= 8'b11111111;
		16'b1010001101110001: data <= 8'b11111111;
		16'b1010001110111110: data <= 8'b11111111;
		16'b1010001110111111: data <= 8'b11111111;
		16'b1010001111000000: data <= 8'b11111111;
		16'b1010001111000001: data <= 8'b11111111;
		16'b1010010001011110: data <= 8'b11111111;
		16'b1010010001011111: data <= 8'b11111111;
		16'b1010010001100000: data <= 8'b11111111;
		16'b1010010001100001: data <= 8'b11111111;
		16'b1010010010101110: data <= 8'b11111111;
		16'b1010010010101111: data <= 8'b11111111;
		16'b1010010010110000: data <= 8'b11111111;
		16'b1010010010110001: data <= 8'b11111111;
		16'b1010010101001110: data <= 8'b11111111;
		16'b1010010101001111: data <= 8'b11111111;
		16'b1010010101010000: data <= 8'b11111111;
		16'b1010010101010001: data <= 8'b11111111;
		16'b1010010110011110: data <= 8'b11111111;
		16'b1010010110011111: data <= 8'b11111111;
		16'b1010010110100000: data <= 8'b11111111;
		16'b1010010110100001: data <= 8'b11111111;
		16'b1010011000111110: data <= 8'b11111111;
		16'b1010011000111111: data <= 8'b11111111;
		16'b1010011001000000: data <= 8'b11111111;
		16'b1010011001000001: data <= 8'b11111111;
		16'b1010011010001110: data <= 8'b11111111;
		16'b1010011010001111: data <= 8'b11111111;
		16'b1010011010010000: data <= 8'b11111111;
		16'b1010011010010001: data <= 8'b11111111;
		16'b1010011100101110: data <= 8'b11111111;
		16'b1010011100101111: data <= 8'b11111111;
		16'b1010011100110000: data <= 8'b11111111;
		16'b1010011100110001: data <= 8'b11111111;
		16'b1010011101111110: data <= 8'b11111111;
		16'b1010011101111111: data <= 8'b11111111;
		16'b1010011110000000: data <= 8'b11111111;
		16'b1010011110000001: data <= 8'b11111111;
		16'b1010100000011110: data <= 8'b11111111;
		16'b1010100000011111: data <= 8'b11111111;
		16'b1010100000100000: data <= 8'b11111111;
		16'b1010100000100001: data <= 8'b11111111;
		16'b1010100001101110: data <= 8'b11111111;
		16'b1010100001101111: data <= 8'b11111111;
		16'b1010100001110000: data <= 8'b11111111;
		16'b1010100001110001: data <= 8'b11111111;
		16'b1010100100001110: data <= 8'b11111111;
		16'b1010100100001111: data <= 8'b11111111;
		16'b1010100100010000: data <= 8'b11111111;
		16'b1010100100010001: data <= 8'b11111111;
		16'b1010100101011110: data <= 8'b11111111;
		16'b1010100101011111: data <= 8'b11111111;
		16'b1010100101100000: data <= 8'b11111111;
		16'b1010100101100001: data <= 8'b11111111;
		16'b1010100111111110: data <= 8'b11111111;
		16'b1010100111111111: data <= 8'b11111111;
		16'b1010101000000000: data <= 8'b11111111;
		16'b1010101000000001: data <= 8'b11111111;
		16'b1010101001001110: data <= 8'b11111111;
		16'b1010101001001111: data <= 8'b11111111;
		16'b1010101001010000: data <= 8'b11111111;
		16'b1010101001010001: data <= 8'b11111111;
		16'b1010101011101110: data <= 8'b11111111;
		16'b1010101011101111: data <= 8'b11111111;
		16'b1010101011110000: data <= 8'b11111111;
		16'b1010101011110001: data <= 8'b11111111;
		16'b1010101100111110: data <= 8'b11111111;
		16'b1010101100111111: data <= 8'b11111111;
		16'b1010101101000000: data <= 8'b11111111;
		16'b1010101101000001: data <= 8'b11111111;
		16'b1010101111011110: data <= 8'b11111111;
		16'b1010101111011111: data <= 8'b11111111;
		16'b1010101111100000: data <= 8'b11111111;
		16'b1010101111100001: data <= 8'b11111111;
		16'b1010110000101110: data <= 8'b11111111;
		16'b1010110000101111: data <= 8'b11111111;
		16'b1010110000110000: data <= 8'b11111111;
		16'b1010110000110001: data <= 8'b11111111;
		16'b1010110011001110: data <= 8'b11111111;
		16'b1010110011001111: data <= 8'b11111111;
		16'b1010110011010000: data <= 8'b11111111;
		16'b1010110011010001: data <= 8'b11111111;
		16'b1010110100011110: data <= 8'b11111111;
		16'b1010110100011111: data <= 8'b11111111;
		16'b1010110100100000: data <= 8'b11111111;
		16'b1010110100100001: data <= 8'b11111111;
		16'b1010110110111110: data <= 8'b11111111;
		16'b1010110110111111: data <= 8'b11111111;
		16'b1010110111000000: data <= 8'b11111111;
		16'b1010110111000001: data <= 8'b11111111;
		16'b1010111000001110: data <= 8'b11111111;
		16'b1010111000001111: data <= 8'b11111111;
		16'b1010111000010000: data <= 8'b11111111;
		16'b1010111000010001: data <= 8'b11111111;
		16'b1010111010101110: data <= 8'b11111111;
		16'b1010111010101111: data <= 8'b11111111;
		16'b1010111010110000: data <= 8'b11111111;
		16'b1010111010110001: data <= 8'b11111111;
		16'b1010111011111110: data <= 8'b11111111;
		16'b1010111011111111: data <= 8'b11111111;
		16'b1010111100000000: data <= 8'b11111111;
		16'b1010111100000001: data <= 8'b11111111;
		16'b1010111110011110: data <= 8'b11111111;
		16'b1010111110011111: data <= 8'b11111111;
		16'b1010111110100000: data <= 8'b11111111;
		16'b1010111110100001: data <= 8'b11111111;
		16'b1010111111101110: data <= 8'b11111111;
		16'b1010111111101111: data <= 8'b11111111;
		16'b1010111111110000: data <= 8'b11111111;
		16'b1010111111110001: data <= 8'b11111111;
		16'b1011000010001110: data <= 8'b11111111;
		16'b1011000010001111: data <= 8'b11111111;
		16'b1011000010010000: data <= 8'b11111111;
		16'b1011000010010001: data <= 8'b11111111;
		16'b1011000011011110: data <= 8'b11111111;
		16'b1011000011011111: data <= 8'b11111111;
		16'b1011000011100000: data <= 8'b11111111;
		16'b1011000011100001: data <= 8'b11111111;
		16'b1011000101111110: data <= 8'b11111111;
		16'b1011000101111111: data <= 8'b11111111;
		16'b1011000110000000: data <= 8'b11111111;
		16'b1011000110000001: data <= 8'b11111111;
		16'b1011000111001110: data <= 8'b11111111;
		16'b1011000111001111: data <= 8'b11111111;
		16'b1011000111010000: data <= 8'b11111111;
		16'b1011000111010001: data <= 8'b11111111;
		16'b1011001001101110: data <= 8'b11111111;
		16'b1011001001101111: data <= 8'b11111111;
		16'b1011001001110000: data <= 8'b11111111;
		16'b1011001001110001: data <= 8'b11111111;
		16'b1011001010111110: data <= 8'b11111111;
		16'b1011001010111111: data <= 8'b11111111;
		16'b1011001011000000: data <= 8'b11111111;
		16'b1011001011000001: data <= 8'b11111111;
		16'b1011001101011110: data <= 8'b11111111;
		16'b1011001101011111: data <= 8'b11111111;
		16'b1011001101100000: data <= 8'b11111111;
		16'b1011001101100001: data <= 8'b11111111;
		16'b1011001110101110: data <= 8'b11111111;
		16'b1011001110101111: data <= 8'b11111111;
		16'b1011001110110000: data <= 8'b11111111;
		16'b1011001110110001: data <= 8'b11111111;
		16'b1011010001001110: data <= 8'b11111111;
		16'b1011010001001111: data <= 8'b11111111;
		16'b1011010001010000: data <= 8'b11111111;
		16'b1011010001010001: data <= 8'b11111111;
		16'b1011010010011110: data <= 8'b11111111;
		16'b1011010010011111: data <= 8'b11111111;
		16'b1011010010100000: data <= 8'b11111111;
		16'b1011010010100001: data <= 8'b11111111;
		16'b1011010100111110: data <= 8'b11111111;
		16'b1011010100111111: data <= 8'b11111111;
		16'b1011010101000000: data <= 8'b11111111;
		16'b1011010101000001: data <= 8'b11111111;
		16'b1011010110001110: data <= 8'b11111111;
		16'b1011010110001111: data <= 8'b11111111;
		16'b1011010110010000: data <= 8'b11111111;
		16'b1011010110010001: data <= 8'b11111111;
		16'b1011011000101110: data <= 8'b11111111;
		16'b1011011000101111: data <= 8'b11111111;
		16'b1011011000110000: data <= 8'b11111111;
		16'b1011011000110001: data <= 8'b11111111;
		16'b1011011001111110: data <= 8'b11111111;
		16'b1011011001111111: data <= 8'b11111111;
		16'b1011011010000000: data <= 8'b11111111;
		16'b1011011010000001: data <= 8'b11111111;
		16'b1011011100011110: data <= 8'b11111111;
		16'b1011011100011111: data <= 8'b11111111;
		16'b1011011100100000: data <= 8'b11111111;
		16'b1011011100100001: data <= 8'b11111111;
		16'b1011011101101110: data <= 8'b11111111;
		16'b1011011101101111: data <= 8'b11111111;
		16'b1011011101110000: data <= 8'b11111111;
		16'b1011011101110001: data <= 8'b11111111;
		16'b1011100000001110: data <= 8'b11111111;
		16'b1011100000001111: data <= 8'b11111111;
		16'b1011100000010000: data <= 8'b11111111;
		16'b1011100000010001: data <= 8'b11111111;
		16'b1011100001011110: data <= 8'b11111111;
		16'b1011100001011111: data <= 8'b11111111;
		16'b1011100001100000: data <= 8'b11111111;
		16'b1011100001100001: data <= 8'b11111111;
		16'b1011100011111110: data <= 8'b11111111;
		16'b1011100011111111: data <= 8'b11111111;
		16'b1011100100000000: data <= 8'b11111111;
		16'b1011100100000001: data <= 8'b11111111;
		16'b1011100101001110: data <= 8'b11111111;
		16'b1011100101001111: data <= 8'b11111111;
		16'b1011100101010000: data <= 8'b11111111;
		16'b1011100101010001: data <= 8'b11111111;
		16'b1011100111101110: data <= 8'b11111111;
		16'b1011100111101111: data <= 8'b11111111;
		16'b1011100111110000: data <= 8'b11111111;
		16'b1011100111110001: data <= 8'b11111111;
		16'b1011101000111110: data <= 8'b11111111;
		16'b1011101000111111: data <= 8'b11111111;
		16'b1011101001000000: data <= 8'b11111111;
		16'b1011101001000001: data <= 8'b11111111;
		16'b1011101011011110: data <= 8'b11111111;
		16'b1011101011011111: data <= 8'b11111111;
		16'b1011101011100000: data <= 8'b11111111;
		16'b1011101011100001: data <= 8'b11111111;
		16'b1011101100101110: data <= 8'b11111111;
		16'b1011101100101111: data <= 8'b11111111;
		16'b1011101100110000: data <= 8'b11111111;
		16'b1011101100110001: data <= 8'b11111111;
		16'b1011101111001110: data <= 8'b11111111;
		16'b1011101111001111: data <= 8'b11111111;
		16'b1011101111010000: data <= 8'b11111111;
		16'b1011101111010001: data <= 8'b11111111;
		16'b1011110000011110: data <= 8'b11111111;
		16'b1011110000011111: data <= 8'b11111111;
		16'b1011110000100000: data <= 8'b11111111;
		16'b1011110000100001: data <= 8'b11111111;
		16'b1011110010111110: data <= 8'b11111111;
		16'b1011110010111111: data <= 8'b11111111;
		16'b1011110011000000: data <= 8'b11111111;
		16'b1011110011000001: data <= 8'b11111111;
		16'b1011110100001110: data <= 8'b11111111;
		16'b1011110100001111: data <= 8'b11111111;
		16'b1011110100010000: data <= 8'b11111111;
		16'b1011110100010001: data <= 8'b11111111;
		16'b1011110110101110: data <= 8'b11111111;
		16'b1011110110101111: data <= 8'b11111111;
		16'b1011110110110000: data <= 8'b11111111;
		16'b1011110110110001: data <= 8'b11111111;
		16'b1011110111111110: data <= 8'b11111111;
		16'b1011110111111111: data <= 8'b11111111;
		16'b1011111000000000: data <= 8'b11111111;
		16'b1011111000000001: data <= 8'b11111111;
		16'b1011111010011110: data <= 8'b11111111;
		16'b1011111010011111: data <= 8'b11111111;
		16'b1011111010100000: data <= 8'b11111111;
		16'b1011111010100001: data <= 8'b11111111;
		16'b1011111011101110: data <= 8'b11111111;
		16'b1011111011101111: data <= 8'b11111111;
		16'b1011111011110000: data <= 8'b11111111;
		16'b1011111011110001: data <= 8'b11111111;
		16'b1011111110001110: data <= 8'b11111111;
		16'b1011111110001111: data <= 8'b11111111;
		16'b1011111110010000: data <= 8'b11111111;
		16'b1011111110010001: data <= 8'b11111111;
		16'b1011111111011110: data <= 8'b11111111;
		16'b1011111111011111: data <= 8'b11111111;
		16'b1011111111100000: data <= 8'b11111111;
		16'b1011111111100001: data <= 8'b11111111;
		16'b1100000001111110: data <= 8'b11111111;
		16'b1100000001111111: data <= 8'b11111111;
		16'b1100000010000000: data <= 8'b11111111;
		16'b1100000010000001: data <= 8'b11111111;
		16'b1100000011001110: data <= 8'b11111111;
		16'b1100000011001111: data <= 8'b11111111;
		16'b1100000011010000: data <= 8'b11111111;
		16'b1100000011010001: data <= 8'b11111111;
		16'b1100000101101110: data <= 8'b11111111;
		16'b1100000101101111: data <= 8'b11111111;
		16'b1100000101110000: data <= 8'b11111111;
		16'b1100000101110001: data <= 8'b11111111;
		16'b1100000110111110: data <= 8'b11111111;
		16'b1100000110111111: data <= 8'b11111111;
		16'b1100000111000000: data <= 8'b11111111;
		16'b1100000111000001: data <= 8'b11111111;
		16'b1100001001011110: data <= 8'b11111111;
		16'b1100001001011111: data <= 8'b11111111;
		16'b1100001001100000: data <= 8'b11111111;
		16'b1100001001100001: data <= 8'b11111111;
		16'b1100001010101110: data <= 8'b11111111;
		16'b1100001010101111: data <= 8'b11111111;
		16'b1100001010110000: data <= 8'b11111111;
		16'b1100001010110001: data <= 8'b11111111;
		16'b1100001101001110: data <= 8'b11111111;
		16'b1100001101001111: data <= 8'b11111111;
		16'b1100001101010000: data <= 8'b11111111;
		16'b1100001101010001: data <= 8'b11111111;
		16'b1100001110011110: data <= 8'b11111111;
		16'b1100001110011111: data <= 8'b11111111;
		16'b1100001110100000: data <= 8'b11111111;
		16'b1100001110100001: data <= 8'b11111111;
		16'b1100010000111110: data <= 8'b11111111;
		16'b1100010000111111: data <= 8'b11111111;
		16'b1100010001000000: data <= 8'b11111111;
		16'b1100010001000001: data <= 8'b11111111;
		16'b1100010010001110: data <= 8'b11111111;
		16'b1100010010001111: data <= 8'b11111111;
		16'b1100010010010000: data <= 8'b11111111;
		16'b1100010010010001: data <= 8'b11111111;
		16'b1100010100101110: data <= 8'b11111111;
		16'b1100010100101111: data <= 8'b11111111;
		16'b1100010100110000: data <= 8'b11111111;
		16'b1100010100110001: data <= 8'b11111111;
		16'b1100010101111110: data <= 8'b11111111;
		16'b1100010101111111: data <= 8'b11111111;
		16'b1100010110000000: data <= 8'b11111111;
		16'b1100010110000001: data <= 8'b11111111;
		16'b1100011000011110: data <= 8'b11111111;
		16'b1100011000011111: data <= 8'b11111111;
		16'b1100011000100000: data <= 8'b11111111;
		16'b1100011000100001: data <= 8'b11111111;
		16'b1100011001101110: data <= 8'b11111111;
		16'b1100011001101111: data <= 8'b11111111;
		16'b1100011001110000: data <= 8'b11111111;
		16'b1100011001110001: data <= 8'b11111111;
		16'b1100011100001110: data <= 8'b11111111;
		16'b1100011100001111: data <= 8'b11111111;
		16'b1100011100010000: data <= 8'b11111111;
		16'b1100011100010001: data <= 8'b11111111;
		16'b1100011101011110: data <= 8'b11111111;
		16'b1100011101011111: data <= 8'b11111111;
		16'b1100011101100000: data <= 8'b11111111;
		16'b1100011101100001: data <= 8'b11111111;
		16'b1100011111111110: data <= 8'b11111111;
		16'b1100011111111111: data <= 8'b11111111;
		16'b1100100000000000: data <= 8'b11111111;
		16'b1100100000000001: data <= 8'b11111111;
		16'b1100100001001110: data <= 8'b11111111;
		16'b1100100001001111: data <= 8'b11111111;
		16'b1100100001010000: data <= 8'b11111111;
		16'b1100100001010001: data <= 8'b11111111;
		16'b1100100011101110: data <= 8'b11111111;
		16'b1100100011101111: data <= 8'b11111111;
		16'b1100100011110000: data <= 8'b11111111;
		16'b1100100011110001: data <= 8'b11111111;
		16'b1100100100111110: data <= 8'b11111111;
		16'b1100100100111111: data <= 8'b11111111;
		16'b1100100101000000: data <= 8'b11111111;
		16'b1100100101000001: data <= 8'b11111111;
		16'b1100100111011110: data <= 8'b11111111;
		16'b1100100111011111: data <= 8'b11111111;
		16'b1100100111100000: data <= 8'b11111111;
		16'b1100100111100001: data <= 8'b11111111;
		16'b1100101000101110: data <= 8'b11111111;
		16'b1100101000101111: data <= 8'b11111111;
		16'b1100101000110000: data <= 8'b11111111;
		16'b1100101000110001: data <= 8'b11111111;
		16'b1100101011001110: data <= 8'b11111111;
		16'b1100101011001111: data <= 8'b11111111;
		16'b1100101011010000: data <= 8'b11111111;
		16'b1100101011010001: data <= 8'b11111111;
		16'b1100101100011110: data <= 8'b11111111;
		16'b1100101100011111: data <= 8'b11111111;
		16'b1100101100100000: data <= 8'b11111111;
		16'b1100101100100001: data <= 8'b11111111;
		16'b1100101110111110: data <= 8'b11111111;
		16'b1100101110111111: data <= 8'b11111111;
		16'b1100101111000000: data <= 8'b11111111;
		16'b1100101111000001: data <= 8'b11111111;
		16'b1100110000001110: data <= 8'b11111111;
		16'b1100110000001111: data <= 8'b11111111;
		16'b1100110000010000: data <= 8'b11111111;
		16'b1100110000010001: data <= 8'b11111111;
		16'b1100110010101110: data <= 8'b11111111;
		16'b1100110010101111: data <= 8'b11111111;
		16'b1100110010110000: data <= 8'b11111111;
		16'b1100110010110001: data <= 8'b11111111;
		16'b1100110011111110: data <= 8'b11111111;
		16'b1100110011111111: data <= 8'b11111111;
		16'b1100110100000000: data <= 8'b11111111;
		16'b1100110100000001: data <= 8'b11111111;
		16'b1100110110011110: data <= 8'b11111111;
		16'b1100110110011111: data <= 8'b11111111;
		16'b1100110110100000: data <= 8'b11111111;
		16'b1100110110100001: data <= 8'b11111111;
		16'b1100110111101110: data <= 8'b11111111;
		16'b1100110111101111: data <= 8'b11111111;
		16'b1100110111110000: data <= 8'b11111111;
		16'b1100110111110001: data <= 8'b11111111;
		16'b1100111010001110: data <= 8'b11111111;
		16'b1100111010001111: data <= 8'b11111111;
		16'b1100111010010000: data <= 8'b11111111;
		16'b1100111010010001: data <= 8'b11111111;
		16'b1100111011011110: data <= 8'b11111111;
		16'b1100111011011111: data <= 8'b11111111;
		16'b1100111011100000: data <= 8'b11111111;
		16'b1100111011100001: data <= 8'b11111111;
		16'b1100111101111110: data <= 8'b11111111;
		16'b1100111101111111: data <= 8'b11111111;
		16'b1100111110000000: data <= 8'b11111111;
		16'b1100111110000001: data <= 8'b11111111;
		16'b1100111111001110: data <= 8'b11111111;
		16'b1100111111001111: data <= 8'b11111111;
		16'b1100111111010000: data <= 8'b11111111;
		16'b1100111111010001: data <= 8'b11111111;
		16'b1101000001101110: data <= 8'b11111111;
		16'b1101000001101111: data <= 8'b11111111;
		16'b1101000001110000: data <= 8'b11111111;
		16'b1101000001110001: data <= 8'b11111111;
		16'b1101000010111110: data <= 8'b11111111;
		16'b1101000010111111: data <= 8'b11111111;
		16'b1101000011000000: data <= 8'b11111111;
		16'b1101000011000001: data <= 8'b11111111;
		16'b1101000101011110: data <= 8'b11111111;
		16'b1101000101011111: data <= 8'b11111111;
		16'b1101000101100000: data <= 8'b11111111;
		16'b1101000101100001: data <= 8'b11111111;
		16'b1101000110101110: data <= 8'b11111111;
		16'b1101000110101111: data <= 8'b11111111;
		16'b1101000110110000: data <= 8'b11111111;
		16'b1101000110110001: data <= 8'b11111111;
		16'b1101001001001110: data <= 8'b11111111;
		16'b1101001001001111: data <= 8'b11111111;
		16'b1101001001010000: data <= 8'b11111111;
		16'b1101001001010001: data <= 8'b11111111;
		16'b1101001010011110: data <= 8'b11111111;
		16'b1101001010011111: data <= 8'b11111111;
		16'b1101001010100000: data <= 8'b11111111;
		16'b1101001010100001: data <= 8'b11111111;
		16'b1101001100111110: data <= 8'b11111111;
		16'b1101001100111111: data <= 8'b11111111;
		16'b1101001101000000: data <= 8'b11111111;
		16'b1101001101000001: data <= 8'b11111111;
		16'b1101001110001110: data <= 8'b11111111;
		16'b1101001110001111: data <= 8'b11111111;
		16'b1101001110010000: data <= 8'b11111111;
		16'b1101001110010001: data <= 8'b11111111;
		16'b1101010000101110: data <= 8'b11111111;
		16'b1101010000101111: data <= 8'b11111111;
		16'b1101010000110000: data <= 8'b11111111;
		16'b1101010000110001: data <= 8'b11111111;
		16'b1101010001111110: data <= 8'b11111111;
		16'b1101010001111111: data <= 8'b11111111;
		16'b1101010010000000: data <= 8'b11111111;
		16'b1101010010000001: data <= 8'b11111111;
		16'b1101010100011110: data <= 8'b11111111;
		16'b1101010100011111: data <= 8'b11111111;
		16'b1101010100100000: data <= 8'b11111111;
		16'b1101010100100001: data <= 8'b11111111;
		16'b1101010101101110: data <= 8'b11111111;
		16'b1101010101101111: data <= 8'b11111111;
		16'b1101010101110000: data <= 8'b11111111;
		16'b1101010101110001: data <= 8'b11111111;
		16'b1101011000001110: data <= 8'b11111111;
		16'b1101011000001111: data <= 8'b11111111;
		16'b1101011000010000: data <= 8'b11111111;
		16'b1101011000010001: data <= 8'b11111111;
		16'b1101011001011110: data <= 8'b11111111;
		16'b1101011001011111: data <= 8'b11111111;
		16'b1101011001100000: data <= 8'b11111111;
		16'b1101011001100001: data <= 8'b11111111;
		16'b1101011011111110: data <= 8'b11111111;
		16'b1101011011111111: data <= 8'b11111111;
		16'b1101011100000000: data <= 8'b11111111;
		16'b1101011100000001: data <= 8'b11111111;
		16'b1101011101001110: data <= 8'b11111111;
		16'b1101011101001111: data <= 8'b11111111;
		16'b1101011101010000: data <= 8'b11111111;
		16'b1101011101010001: data <= 8'b11111111;
		16'b1101011111101110: data <= 8'b11111111;
		16'b1101011111101111: data <= 8'b11111111;
		16'b1101011111110000: data <= 8'b11111111;
		16'b1101011111110001: data <= 8'b11111111;
		16'b1101100000111110: data <= 8'b11111111;
		16'b1101100000111111: data <= 8'b11111111;
		16'b1101100001000000: data <= 8'b11111111;
		16'b1101100001000001: data <= 8'b11111111;
		16'b1101100011011110: data <= 8'b11111111;
		16'b1101100011011111: data <= 8'b11111111;
		16'b1101100011100000: data <= 8'b11111111;
		16'b1101100011100001: data <= 8'b11111111;
		16'b1101100100101110: data <= 8'b11111111;
		16'b1101100100101111: data <= 8'b11111111;
		16'b1101100100110000: data <= 8'b11111111;
		16'b1101100100110001: data <= 8'b11111111;
		16'b1101100111001110: data <= 8'b11111111;
		16'b1101100111001111: data <= 8'b11111111;
		16'b1101100111010000: data <= 8'b11111111;
		16'b1101100111010001: data <= 8'b11111111;
		16'b1101101000011110: data <= 8'b11111111;
		16'b1101101000011111: data <= 8'b11111111;
		16'b1101101000100000: data <= 8'b11111111;
		16'b1101101000100001: data <= 8'b11111111;
		16'b1101101010111110: data <= 8'b11111111;
		16'b1101101010111111: data <= 8'b11111111;
		16'b1101101011000000: data <= 8'b11111111;
		16'b1101101011000001: data <= 8'b11111111;
		16'b1101101100001110: data <= 8'b11111111;
		16'b1101101100001111: data <= 8'b11111111;
		16'b1101101100010000: data <= 8'b11111111;
		16'b1101101100010001: data <= 8'b11111111;
		16'b1101101110101110: data <= 8'b11111111;
		16'b1101101110101111: data <= 8'b11111111;
		16'b1101101110110000: data <= 8'b11111111;
		16'b1101101110110001: data <= 8'b11111111;
		16'b1101101111111110: data <= 8'b11111111;
		16'b1101101111111111: data <= 8'b11111111;
		16'b1101110000000000: data <= 8'b11111111;
		16'b1101110000000001: data <= 8'b11111111;
		16'b1101110010011110: data <= 8'b11111111;
		16'b1101110010011111: data <= 8'b11111111;
		16'b1101110010100000: data <= 8'b11111111;
		16'b1101110010100001: data <= 8'b11111111;
		16'b1101110011101110: data <= 8'b11111111;
		16'b1101110011101111: data <= 8'b11111111;
		16'b1101110011110000: data <= 8'b11111111;
		16'b1101110011110001: data <= 8'b11111111;
		16'b1101110110001110: data <= 8'b11111111;
		16'b1101110110001111: data <= 8'b11111111;
		16'b1101110110010000: data <= 8'b11111111;
		16'b1101110110010001: data <= 8'b11111111;
		16'b1101110111011110: data <= 8'b11111111;
		16'b1101110111011111: data <= 8'b11111111;
		16'b1101110111100000: data <= 8'b11111111;
		16'b1101110111100001: data <= 8'b11111111;
		16'b1101111001111110: data <= 8'b11111111;
		16'b1101111001111111: data <= 8'b11111111;
		16'b1101111010000000: data <= 8'b11111111;
		16'b1101111010000001: data <= 8'b11111111;
		16'b1101111011001110: data <= 8'b11111111;
		16'b1101111011001111: data <= 8'b11111111;
		16'b1101111011010000: data <= 8'b11111111;
		16'b1101111011010001: data <= 8'b11111111;
		16'b1101111101101110: data <= 8'b11111111;
		16'b1101111101101111: data <= 8'b11111111;
		16'b1101111101110000: data <= 8'b11111111;
		16'b1101111101110001: data <= 8'b11111111;
		16'b1101111110111110: data <= 8'b11111111;
		16'b1101111110111111: data <= 8'b11111111;
		16'b1101111111000000: data <= 8'b11111111;
		16'b1101111111000001: data <= 8'b11111111;
		16'b1110000001011110: data <= 8'b11111111;
		16'b1110000001011111: data <= 8'b11111111;
		16'b1110000001100000: data <= 8'b11111111;
		16'b1110000001100001: data <= 8'b11111111;
		16'b1110000010101110: data <= 8'b11111111;
		16'b1110000010101111: data <= 8'b11111111;
		16'b1110000010110000: data <= 8'b11111111;
		16'b1110000010110001: data <= 8'b11111111;
		default: data <= 8'b00000000;
	endcase
end

endmodule
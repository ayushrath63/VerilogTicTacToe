module score_rom(
//inputs
clk, addr, 
//outputs
data);

(* rom_style = "block" *)

input wire clk;
input wire [9:0] addr;
output reg [7:0] data;

reg [9:0] addr_reg;

always @ (posedge clk)
	addr_reg <= addr;

always @ (*)
begin
	case(addr)
		10'b0000000000: data <= 8'b11111111;
		10'b0000000001: data <= 8'b11111111;
		10'b0000000010: data <= 8'b11111111;
		10'b0000000100: data <= 8'b11111111;
		10'b0000001001: data <= 8'b11111111;
		10'b0000001010: data <= 8'b11111111;
		10'b0000001101: data <= 8'b11111111;
		10'b0000010001: data <= 8'b11111111;
		10'b0000010011: data <= 8'b11111111;
		10'b0000010100: data <= 8'b11111111;
		10'b0000010101: data <= 8'b11111111;
		10'b0000010111: data <= 8'b11111111;
		10'b0000011000: data <= 8'b11111111;
		10'b0000011101: data <= 8'b11111111;
		10'b0000100001: data <= 8'b11111111;
		10'b0000100011: data <= 8'b11111111;
		10'b0000100101: data <= 8'b11111111;
		10'b0000101001: data <= 8'b11111111;
		10'b0000101100: data <= 8'b11111111;
		10'b0000101111: data <= 8'b11111111;
		10'b0000110001: data <= 8'b11111111;
		10'b0000110100: data <= 8'b11111111;
		10'b0000111000: data <= 8'b11111111;
		10'b0000111010: data <= 8'b11111111;
		10'b0000111101: data <= 8'b11111111;
		10'b0000111110: data <= 8'b11111111;
		10'b0001000001: data <= 8'b11111111;
		10'b0001000010: data <= 8'b11111111;
		10'b0001000011: data <= 8'b11111111;
		10'b0001000100: data <= 8'b11111111;
		10'b0001000110: data <= 8'b11111111;
		10'b0001001010: data <= 8'b11111111;
		10'b0001001011: data <= 8'b11111111;
		10'b0001001100: data <= 8'b11111111;
		10'b0001001101: data <= 8'b11111111;
		10'b0001010001: data <= 8'b11111111;
		10'b0001010101: data <= 8'b11111111;
		10'b0001010110: data <= 8'b11111111;
		10'b0001010111: data <= 8'b11111111;
		10'b0001011001: data <= 8'b11111111;
		10'b0001011010: data <= 8'b11111111;
		10'b0001011111: data <= 8'b11111111;
		10'b0001100011: data <= 8'b11111111;
		10'b0001100111: data <= 8'b11111111;
		10'b0001101011: data <= 8'b11111111;
		10'b0001101110: data <= 8'b11111111;
		10'b0001110010: data <= 8'b11111111;
		10'b0001110110: data <= 8'b11111111;
		10'b0001111010: data <= 8'b11111111;
		10'b0001111100: data <= 8'b11111111;
		10'b0010000000: data <= 8'b11111111;
		10'b0010000011: data <= 8'b11111111;
		10'b0010000100: data <= 8'b11111111;
		10'b0010001000: data <= 8'b11111111;
		10'b0010001001: data <= 8'b11111111;
		10'b0010001010: data <= 8'b11111111;
		10'b0010001100: data <= 8'b11111111;
		10'b0010001111: data <= 8'b11111111;
		10'b0010010011: data <= 8'b11111111;
		10'b0010010111: data <= 8'b11111111;
		10'b0010011000: data <= 8'b11111111;
		10'b0010011001: data <= 8'b11111111;
		10'b0010011011: data <= 8'b11111111;
		10'b0010011101: data <= 8'b11111111;
		10'b0010100000: data <= 8'b11111111;
		10'b0010100001: data <= 8'b11111111;
		10'b0010100010: data <= 8'b11111111;
		10'b0011000110: data <= 8'b11111111;
		10'b0011000111: data <= 8'b11111111;
		10'b0011001000: data <= 8'b11111111;
		10'b0011001010: data <= 8'b11111111;
		10'b0011001111: data <= 8'b11111111;
		10'b0011010000: data <= 8'b11111111;
		10'b0011010011: data <= 8'b11111111;
		10'b0011010111: data <= 8'b11111111;
		10'b0011011001: data <= 8'b11111111;
		10'b0011011010: data <= 8'b11111111;
		10'b0011011011: data <= 8'b11111111;
		10'b0011011101: data <= 8'b11111111;
		10'b0011011110: data <= 8'b11111111;
		10'b0011100011: data <= 8'b11111111;
		10'b0011100111: data <= 8'b11111111;
		10'b0011101001: data <= 8'b11111111;
		10'b0011101011: data <= 8'b11111111;
		10'b0011101111: data <= 8'b11111111;
		10'b0011110010: data <= 8'b11111111;
		10'b0011110101: data <= 8'b11111111;
		10'b0011110111: data <= 8'b11111111;
		10'b0011111010: data <= 8'b11111111;
		10'b0011111110: data <= 8'b11111111;
		10'b0100000000: data <= 8'b11111111;
		10'b0100000011: data <= 8'b11111111;
		10'b0100000101: data <= 8'b11111111;
		10'b0100000111: data <= 8'b11111111;
		10'b0100001000: data <= 8'b11111111;
		10'b0100001001: data <= 8'b11111111;
		10'b0100001010: data <= 8'b11111111;
		10'b0100001100: data <= 8'b11111111;
		10'b0100010000: data <= 8'b11111111;
		10'b0100010001: data <= 8'b11111111;
		10'b0100010010: data <= 8'b11111111;
		10'b0100010011: data <= 8'b11111111;
		10'b0100010111: data <= 8'b11111111;
		10'b0100011011: data <= 8'b11111111;
		10'b0100011100: data <= 8'b11111111;
		10'b0100011101: data <= 8'b11111111;
		10'b0100011111: data <= 8'b11111111;
		10'b0100100000: data <= 8'b11111111;
		10'b0100100110: data <= 8'b11111111;
		10'b0100101001: data <= 8'b11111111;
		10'b0100101101: data <= 8'b11111111;
		10'b0100110001: data <= 8'b11111111;
		10'b0100110100: data <= 8'b11111111;
		10'b0100111000: data <= 8'b11111111;
		10'b0100111100: data <= 8'b11111111;
		10'b0101000000: data <= 8'b11111111;
		10'b0101000010: data <= 8'b11111111;
		10'b0101000110: data <= 8'b11111111;
		10'b0101001001: data <= 8'b11111111;
		10'b0101001010: data <= 8'b11111111;
		10'b0101001110: data <= 8'b11111111;
		10'b0101001111: data <= 8'b11111111;
		10'b0101010000: data <= 8'b11111111;
		10'b0101010010: data <= 8'b11111111;
		10'b0101010101: data <= 8'b11111111;
		10'b0101011001: data <= 8'b11111111;
		10'b0101011101: data <= 8'b11111111;
		10'b0101011110: data <= 8'b11111111;
		10'b0101011111: data <= 8'b11111111;
		10'b0101100001: data <= 8'b11111111;
		10'b0101100011: data <= 8'b11111111;
		10'b0101100110: data <= 8'b11111111;
		10'b0101100111: data <= 8'b11111111;
		10'b0101101000: data <= 8'b11111111;
		10'b0110011100: data <= 8'b11111111;
		10'b0110011101: data <= 8'b11111111;
		10'b0110011110: data <= 8'b11111111;
		10'b0110100000: data <= 8'b11111111;
		10'b0110100001: data <= 8'b11111111;
		10'b0110100010: data <= 8'b11111111;
		10'b0110100100: data <= 8'b11111111;
		10'b0110100101: data <= 8'b11111111;
		10'b0110100110: data <= 8'b11111111;
		10'b0110101001: data <= 8'b11111111;
		10'b0110101010: data <= 8'b11111111;
		10'b0110111110: data <= 8'b11111111;
		10'b0111000010: data <= 8'b11111111;
		10'b0111000101: data <= 8'b11111111;
		10'b0111001001: data <= 8'b11111111;
		10'b0111001101: data <= 8'b11111111;
		10'b0111011111: data <= 8'b11111111;
		10'b0111100011: data <= 8'b11111111;
		10'b0111100110: data <= 8'b11111111;
		10'b0111100111: data <= 8'b11111111;
		10'b0111101000: data <= 8'b11111111;
		10'b0111101011: data <= 8'b11111111;
		10'b1000000000: data <= 8'b11111111;
		10'b1000000100: data <= 8'b11111111;
		10'b1000000111: data <= 8'b11111111;
		10'b1000001101: data <= 8'b11111111;
		10'b1000001111: data <= 8'b11111111;
		10'b1000100001: data <= 8'b11111111;
		10'b1000100100: data <= 8'b11111111;
		10'b1000100101: data <= 8'b11111111;
		10'b1000100110: data <= 8'b11111111;
		10'b1000101000: data <= 8'b11111111;
		10'b1000101001: data <= 8'b11111111;
		10'b1000101010: data <= 8'b11111111;
		10'b1000101100: data <= 8'b11111111;
		10'b1000101101: data <= 8'b11111111;
		default: data <= 8'b00000000;
	endcase
end

endmodule
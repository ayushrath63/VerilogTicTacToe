module o_rom(
//inputs
clk, addr, 
//outputs
data);

(* rom_style = "block" *)

input wire clk;
input wire [12:0] addr;
output reg [7:0] data;

reg [12:0] addr_reg;

always @ (posedge clk)
	addr_reg <= addr;

always @ (*)
begin
	case(addr)
		13'b0010001111111: data <= 8'b11111111;
		13'b0010010000000: data <= 8'b11111111;
		13'b0010010000001: data <= 8'b11111111;
		13'b0010010000010: data <= 8'b11111111;
		13'b0010010000011: data <= 8'b11111111;
		13'b0010010000100: data <= 8'b11111111;
		13'b0010010000101: data <= 8'b11111111;
		13'b0010010000110: data <= 8'b11111111;
		13'b0010010000111: data <= 8'b11111111;
		13'b0010010001000: data <= 8'b11111111;
		13'b0010010001001: data <= 8'b11111111;
		13'b0010010001010: data <= 8'b11111111;
		13'b0010010001011: data <= 8'b11111111;
		13'b0010010001100: data <= 8'b11111111;
		13'b0010010001101: data <= 8'b11111111;
		13'b0010010001110: data <= 8'b11111111;
		13'b0010010001111: data <= 8'b11111111;
		13'b0010010010000: data <= 8'b11111111;
		13'b0010011001110: data <= 8'b11111111;
		13'b0010011001111: data <= 8'b11111111;
		13'b0010011010000: data <= 8'b11111111;
		13'b0010011010001: data <= 8'b11111111;
		13'b0010011010010: data <= 8'b11111111;
		13'b0010011010011: data <= 8'b11111111;
		13'b0010011010100: data <= 8'b11111111;
		13'b0010011010101: data <= 8'b11111111;
		13'b0010011010110: data <= 8'b11111111;
		13'b0010011010111: data <= 8'b11111111;
		13'b0010011011000: data <= 8'b11111111;
		13'b0010011011001: data <= 8'b11111111;
		13'b0010011011010: data <= 8'b11111111;
		13'b0010011011011: data <= 8'b11111111;
		13'b0010011011100: data <= 8'b11111111;
		13'b0010011011101: data <= 8'b11111111;
		13'b0010011011110: data <= 8'b11111111;
		13'b0010011011111: data <= 8'b11111111;
		13'b0010011100000: data <= 8'b11111111;
		13'b0010011100001: data <= 8'b11111111;
		13'b0010100011101: data <= 8'b11111111;
		13'b0010100011110: data <= 8'b11111111;
		13'b0010100011111: data <= 8'b11111111;
		13'b0010100100000: data <= 8'b11111111;
		13'b0010100100001: data <= 8'b11111111;
		13'b0010100100010: data <= 8'b11111111;
		13'b0010100100011: data <= 8'b11111111;
		13'b0010100100100: data <= 8'b11111111;
		13'b0010100100101: data <= 8'b11111111;
		13'b0010100100110: data <= 8'b11111111;
		13'b0010100100111: data <= 8'b11111111;
		13'b0010100101000: data <= 8'b11111111;
		13'b0010100101001: data <= 8'b11111111;
		13'b0010100101010: data <= 8'b11111111;
		13'b0010100101011: data <= 8'b11111111;
		13'b0010100101100: data <= 8'b11111111;
		13'b0010100101101: data <= 8'b11111111;
		13'b0010100101110: data <= 8'b11111111;
		13'b0010100101111: data <= 8'b11111111;
		13'b0010100110000: data <= 8'b11111111;
		13'b0010100110001: data <= 8'b11111111;
		13'b0010100110010: data <= 8'b11111111;
		13'b0010101101100: data <= 8'b11111111;
		13'b0010101101101: data <= 8'b11111111;
		13'b0010101101110: data <= 8'b11111111;
		13'b0010101101111: data <= 8'b11111111;
		13'b0010101110000: data <= 8'b11111111;
		13'b0010101110001: data <= 8'b11111111;
		13'b0010101110010: data <= 8'b11111111;
		13'b0010101110011: data <= 8'b11111111;
		13'b0010101110100: data <= 8'b11111111;
		13'b0010101110101: data <= 8'b11111111;
		13'b0010101110110: data <= 8'b11111111;
		13'b0010101110111: data <= 8'b11111111;
		13'b0010101111000: data <= 8'b11111111;
		13'b0010101111001: data <= 8'b11111111;
		13'b0010101111010: data <= 8'b11111111;
		13'b0010101111011: data <= 8'b11111111;
		13'b0010101111100: data <= 8'b11111111;
		13'b0010101111101: data <= 8'b11111111;
		13'b0010101111110: data <= 8'b11111111;
		13'b0010101111111: data <= 8'b11111111;
		13'b0010110000000: data <= 8'b11111111;
		13'b0010110000001: data <= 8'b11111111;
		13'b0010110000010: data <= 8'b11111111;
		13'b0010110000011: data <= 8'b11111111;
		13'b0010110111011: data <= 8'b11111111;
		13'b0010110111100: data <= 8'b11111111;
		13'b0010110111101: data <= 8'b11111111;
		13'b0010110111110: data <= 8'b11111111;
		13'b0010110111111: data <= 8'b11111111;
		13'b0010111010000: data <= 8'b11111111;
		13'b0010111010001: data <= 8'b11111111;
		13'b0010111010010: data <= 8'b11111111;
		13'b0010111010011: data <= 8'b11111111;
		13'b0010111010100: data <= 8'b11111111;
		13'b0011000001010: data <= 8'b11111111;
		13'b0011000001011: data <= 8'b11111111;
		13'b0011000001100: data <= 8'b11111111;
		13'b0011000001101: data <= 8'b11111111;
		13'b0011000001110: data <= 8'b11111111;
		13'b0011000100001: data <= 8'b11111111;
		13'b0011000100010: data <= 8'b11111111;
		13'b0011000100011: data <= 8'b11111111;
		13'b0011000100100: data <= 8'b11111111;
		13'b0011000100101: data <= 8'b11111111;
		13'b0011001011001: data <= 8'b11111111;
		13'b0011001011010: data <= 8'b11111111;
		13'b0011001011011: data <= 8'b11111111;
		13'b0011001011100: data <= 8'b11111111;
		13'b0011001011101: data <= 8'b11111111;
		13'b0011001110010: data <= 8'b11111111;
		13'b0011001110011: data <= 8'b11111111;
		13'b0011001110100: data <= 8'b11111111;
		13'b0011001110101: data <= 8'b11111111;
		13'b0011001110110: data <= 8'b11111111;
		13'b0011010101000: data <= 8'b11111111;
		13'b0011010101001: data <= 8'b11111111;
		13'b0011010101010: data <= 8'b11111111;
		13'b0011010101011: data <= 8'b11111111;
		13'b0011010101100: data <= 8'b11111111;
		13'b0011011000011: data <= 8'b11111111;
		13'b0011011000100: data <= 8'b11111111;
		13'b0011011000101: data <= 8'b11111111;
		13'b0011011000110: data <= 8'b11111111;
		13'b0011011000111: data <= 8'b11111111;
		13'b0011011110111: data <= 8'b11111111;
		13'b0011011111000: data <= 8'b11111111;
		13'b0011011111001: data <= 8'b11111111;
		13'b0011011111010: data <= 8'b11111111;
		13'b0011011111011: data <= 8'b11111111;
		13'b0011100010100: data <= 8'b11111111;
		13'b0011100010101: data <= 8'b11111111;
		13'b0011100010110: data <= 8'b11111111;
		13'b0011100010111: data <= 8'b11111111;
		13'b0011100011000: data <= 8'b11111111;
		13'b0011101000110: data <= 8'b11111111;
		13'b0011101000111: data <= 8'b11111111;
		13'b0011101001000: data <= 8'b11111111;
		13'b0011101001001: data <= 8'b11111111;
		13'b0011101001010: data <= 8'b11111111;
		13'b0011101100101: data <= 8'b11111111;
		13'b0011101100110: data <= 8'b11111111;
		13'b0011101100111: data <= 8'b11111111;
		13'b0011101101000: data <= 8'b11111111;
		13'b0011101101001: data <= 8'b11111111;
		13'b0011110010110: data <= 8'b11111111;
		13'b0011110010111: data <= 8'b11111111;
		13'b0011110011000: data <= 8'b11111111;
		13'b0011110011001: data <= 8'b11111111;
		13'b0011110110110: data <= 8'b11111111;
		13'b0011110110111: data <= 8'b11111111;
		13'b0011110111000: data <= 8'b11111111;
		13'b0011110111001: data <= 8'b11111111;
		13'b0011111100110: data <= 8'b11111111;
		13'b0011111100111: data <= 8'b11111111;
		13'b0011111101000: data <= 8'b11111111;
		13'b0011111101001: data <= 8'b11111111;
		13'b0100000000110: data <= 8'b11111111;
		13'b0100000000111: data <= 8'b11111111;
		13'b0100000001000: data <= 8'b11111111;
		13'b0100000001001: data <= 8'b11111111;
		13'b0100000110110: data <= 8'b11111111;
		13'b0100000110111: data <= 8'b11111111;
		13'b0100000111000: data <= 8'b11111111;
		13'b0100000111001: data <= 8'b11111111;
		13'b0100001010110: data <= 8'b11111111;
		13'b0100001010111: data <= 8'b11111111;
		13'b0100001011000: data <= 8'b11111111;
		13'b0100001011001: data <= 8'b11111111;
		13'b0100010000110: data <= 8'b11111111;
		13'b0100010000111: data <= 8'b11111111;
		13'b0100010001000: data <= 8'b11111111;
		13'b0100010001001: data <= 8'b11111111;
		13'b0100010100110: data <= 8'b11111111;
		13'b0100010100111: data <= 8'b11111111;
		13'b0100010101000: data <= 8'b11111111;
		13'b0100010101001: data <= 8'b11111111;
		13'b0100011010110: data <= 8'b11111111;
		13'b0100011010111: data <= 8'b11111111;
		13'b0100011011000: data <= 8'b11111111;
		13'b0100011011001: data <= 8'b11111111;
		13'b0100011110110: data <= 8'b11111111;
		13'b0100011110111: data <= 8'b11111111;
		13'b0100011111000: data <= 8'b11111111;
		13'b0100011111001: data <= 8'b11111111;
		13'b0100100100110: data <= 8'b11111111;
		13'b0100100100111: data <= 8'b11111111;
		13'b0100100101000: data <= 8'b11111111;
		13'b0100100101001: data <= 8'b11111111;
		13'b0100101000110: data <= 8'b11111111;
		13'b0100101000111: data <= 8'b11111111;
		13'b0100101001000: data <= 8'b11111111;
		13'b0100101001001: data <= 8'b11111111;
		13'b0100101110110: data <= 8'b11111111;
		13'b0100101110111: data <= 8'b11111111;
		13'b0100101111000: data <= 8'b11111111;
		13'b0100101111001: data <= 8'b11111111;
		13'b0100110010110: data <= 8'b11111111;
		13'b0100110010111: data <= 8'b11111111;
		13'b0100110011000: data <= 8'b11111111;
		13'b0100110011001: data <= 8'b11111111;
		13'b0100111000110: data <= 8'b11111111;
		13'b0100111000111: data <= 8'b11111111;
		13'b0100111001000: data <= 8'b11111111;
		13'b0100111001001: data <= 8'b11111111;
		13'b0100111100110: data <= 8'b11111111;
		13'b0100111100111: data <= 8'b11111111;
		13'b0100111101000: data <= 8'b11111111;
		13'b0100111101001: data <= 8'b11111111;
		13'b0101000010110: data <= 8'b11111111;
		13'b0101000010111: data <= 8'b11111111;
		13'b0101000011000: data <= 8'b11111111;
		13'b0101000011001: data <= 8'b11111111;
		13'b0101000110110: data <= 8'b11111111;
		13'b0101000110111: data <= 8'b11111111;
		13'b0101000111000: data <= 8'b11111111;
		13'b0101000111001: data <= 8'b11111111;
		13'b0101001100110: data <= 8'b11111111;
		13'b0101001100111: data <= 8'b11111111;
		13'b0101001101000: data <= 8'b11111111;
		13'b0101001101001: data <= 8'b11111111;
		13'b0101010000110: data <= 8'b11111111;
		13'b0101010000111: data <= 8'b11111111;
		13'b0101010001000: data <= 8'b11111111;
		13'b0101010001001: data <= 8'b11111111;
		13'b0101010110110: data <= 8'b11111111;
		13'b0101010110111: data <= 8'b11111111;
		13'b0101010111000: data <= 8'b11111111;
		13'b0101010111001: data <= 8'b11111111;
		13'b0101011010110: data <= 8'b11111111;
		13'b0101011010111: data <= 8'b11111111;
		13'b0101011011000: data <= 8'b11111111;
		13'b0101011011001: data <= 8'b11111111;
		13'b0101100000110: data <= 8'b11111111;
		13'b0101100000111: data <= 8'b11111111;
		13'b0101100001000: data <= 8'b11111111;
		13'b0101100001001: data <= 8'b11111111;
		13'b0101100100110: data <= 8'b11111111;
		13'b0101100100111: data <= 8'b11111111;
		13'b0101100101000: data <= 8'b11111111;
		13'b0101100101001: data <= 8'b11111111;
		13'b0101101010110: data <= 8'b11111111;
		13'b0101101010111: data <= 8'b11111111;
		13'b0101101011000: data <= 8'b11111111;
		13'b0101101011001: data <= 8'b11111111;
		13'b0101101110110: data <= 8'b11111111;
		13'b0101101110111: data <= 8'b11111111;
		13'b0101101111000: data <= 8'b11111111;
		13'b0101101111001: data <= 8'b11111111;
		13'b0101110100110: data <= 8'b11111111;
		13'b0101110100111: data <= 8'b11111111;
		13'b0101110101000: data <= 8'b11111111;
		13'b0101110101001: data <= 8'b11111111;
		13'b0101111000110: data <= 8'b11111111;
		13'b0101111000111: data <= 8'b11111111;
		13'b0101111001000: data <= 8'b11111111;
		13'b0101111001001: data <= 8'b11111111;
		13'b0101111110110: data <= 8'b11111111;
		13'b0101111110111: data <= 8'b11111111;
		13'b0101111111000: data <= 8'b11111111;
		13'b0101111111001: data <= 8'b11111111;
		13'b0110000010110: data <= 8'b11111111;
		13'b0110000010111: data <= 8'b11111111;
		13'b0110000011000: data <= 8'b11111111;
		13'b0110000011001: data <= 8'b11111111;
		13'b0110001000110: data <= 8'b11111111;
		13'b0110001000111: data <= 8'b11111111;
		13'b0110001001000: data <= 8'b11111111;
		13'b0110001001001: data <= 8'b11111111;
		13'b0110001100110: data <= 8'b11111111;
		13'b0110001100111: data <= 8'b11111111;
		13'b0110001101000: data <= 8'b11111111;
		13'b0110001101001: data <= 8'b11111111;
		13'b0110010010110: data <= 8'b11111111;
		13'b0110010010111: data <= 8'b11111111;
		13'b0110010011000: data <= 8'b11111111;
		13'b0110010011001: data <= 8'b11111111;
		13'b0110010110110: data <= 8'b11111111;
		13'b0110010110111: data <= 8'b11111111;
		13'b0110010111000: data <= 8'b11111111;
		13'b0110010111001: data <= 8'b11111111;
		13'b0110011100110: data <= 8'b11111111;
		13'b0110011100111: data <= 8'b11111111;
		13'b0110011101000: data <= 8'b11111111;
		13'b0110011101001: data <= 8'b11111111;
		13'b0110100000110: data <= 8'b11111111;
		13'b0110100000111: data <= 8'b11111111;
		13'b0110100001000: data <= 8'b11111111;
		13'b0110100001001: data <= 8'b11111111;
		13'b0110100110110: data <= 8'b11111111;
		13'b0110100110111: data <= 8'b11111111;
		13'b0110100111000: data <= 8'b11111111;
		13'b0110100111001: data <= 8'b11111111;
		13'b0110101010110: data <= 8'b11111111;
		13'b0110101010111: data <= 8'b11111111;
		13'b0110101011000: data <= 8'b11111111;
		13'b0110101011001: data <= 8'b11111111;
		13'b0110110000110: data <= 8'b11111111;
		13'b0110110000111: data <= 8'b11111111;
		13'b0110110001000: data <= 8'b11111111;
		13'b0110110001001: data <= 8'b11111111;
		13'b0110110100110: data <= 8'b11111111;
		13'b0110110100111: data <= 8'b11111111;
		13'b0110110101000: data <= 8'b11111111;
		13'b0110110101001: data <= 8'b11111111;
		13'b0110111010110: data <= 8'b11111111;
		13'b0110111010111: data <= 8'b11111111;
		13'b0110111011000: data <= 8'b11111111;
		13'b0110111011001: data <= 8'b11111111;
		13'b0110111110110: data <= 8'b11111111;
		13'b0110111110111: data <= 8'b11111111;
		13'b0110111111000: data <= 8'b11111111;
		13'b0110111111001: data <= 8'b11111111;
		13'b0111000100110: data <= 8'b11111111;
		13'b0111000100111: data <= 8'b11111111;
		13'b0111000101000: data <= 8'b11111111;
		13'b0111000101001: data <= 8'b11111111;
		13'b0111001000110: data <= 8'b11111111;
		13'b0111001000111: data <= 8'b11111111;
		13'b0111001001000: data <= 8'b11111111;
		13'b0111001001001: data <= 8'b11111111;
		13'b0111001110110: data <= 8'b11111111;
		13'b0111001110111: data <= 8'b11111111;
		13'b0111001111000: data <= 8'b11111111;
		13'b0111001111001: data <= 8'b11111111;
		13'b0111010010110: data <= 8'b11111111;
		13'b0111010010111: data <= 8'b11111111;
		13'b0111010011000: data <= 8'b11111111;
		13'b0111010011001: data <= 8'b11111111;
		13'b0111011000110: data <= 8'b11111111;
		13'b0111011000111: data <= 8'b11111111;
		13'b0111011001000: data <= 8'b11111111;
		13'b0111011001001: data <= 8'b11111111;
		13'b0111011100110: data <= 8'b11111111;
		13'b0111011100111: data <= 8'b11111111;
		13'b0111011101000: data <= 8'b11111111;
		13'b0111011101001: data <= 8'b11111111;
		13'b0111100010110: data <= 8'b11111111;
		13'b0111100010111: data <= 8'b11111111;
		13'b0111100011000: data <= 8'b11111111;
		13'b0111100011001: data <= 8'b11111111;
		13'b0111100110110: data <= 8'b11111111;
		13'b0111100110111: data <= 8'b11111111;
		13'b0111100111000: data <= 8'b11111111;
		13'b0111100111001: data <= 8'b11111111;
		13'b0111101100110: data <= 8'b11111111;
		13'b0111101100111: data <= 8'b11111111;
		13'b0111101101000: data <= 8'b11111111;
		13'b0111101101001: data <= 8'b11111111;
		13'b0111110000110: data <= 8'b11111111;
		13'b0111110000111: data <= 8'b11111111;
		13'b0111110001000: data <= 8'b11111111;
		13'b0111110001001: data <= 8'b11111111;
		13'b0111110110110: data <= 8'b11111111;
		13'b0111110110111: data <= 8'b11111111;
		13'b0111110111000: data <= 8'b11111111;
		13'b0111110111001: data <= 8'b11111111;
		13'b0111111010110: data <= 8'b11111111;
		13'b0111111010111: data <= 8'b11111111;
		13'b0111111011000: data <= 8'b11111111;
		13'b0111111011001: data <= 8'b11111111;
		13'b1000000000110: data <= 8'b11111111;
		13'b1000000000111: data <= 8'b11111111;
		13'b1000000001000: data <= 8'b11111111;
		13'b1000000001001: data <= 8'b11111111;
		13'b1000000100110: data <= 8'b11111111;
		13'b1000000100111: data <= 8'b11111111;
		13'b1000000101000: data <= 8'b11111111;
		13'b1000000101001: data <= 8'b11111111;
		13'b1000001010110: data <= 8'b11111111;
		13'b1000001010111: data <= 8'b11111111;
		13'b1000001011000: data <= 8'b11111111;
		13'b1000001011001: data <= 8'b11111111;
		13'b1000001110110: data <= 8'b11111111;
		13'b1000001110111: data <= 8'b11111111;
		13'b1000001111000: data <= 8'b11111111;
		13'b1000001111001: data <= 8'b11111111;
		13'b1000010100110: data <= 8'b11111111;
		13'b1000010100111: data <= 8'b11111111;
		13'b1000010101000: data <= 8'b11111111;
		13'b1000010101001: data <= 8'b11111111;
		13'b1000011000110: data <= 8'b11111111;
		13'b1000011000111: data <= 8'b11111111;
		13'b1000011001000: data <= 8'b11111111;
		13'b1000011001001: data <= 8'b11111111;
		13'b1000011110110: data <= 8'b11111111;
		13'b1000011110111: data <= 8'b11111111;
		13'b1000011111000: data <= 8'b11111111;
		13'b1000011111001: data <= 8'b11111111;
		13'b1000100010110: data <= 8'b11111111;
		13'b1000100010111: data <= 8'b11111111;
		13'b1000100011000: data <= 8'b11111111;
		13'b1000100011001: data <= 8'b11111111;
		13'b1000101000110: data <= 8'b11111111;
		13'b1000101000111: data <= 8'b11111111;
		13'b1000101001000: data <= 8'b11111111;
		13'b1000101001001: data <= 8'b11111111;
		13'b1000101100110: data <= 8'b11111111;
		13'b1000101100111: data <= 8'b11111111;
		13'b1000101101000: data <= 8'b11111111;
		13'b1000101101001: data <= 8'b11111111;
		13'b1000110010110: data <= 8'b11111111;
		13'b1000110010111: data <= 8'b11111111;
		13'b1000110011000: data <= 8'b11111111;
		13'b1000110011001: data <= 8'b11111111;
		13'b1000110011010: data <= 8'b11111111;
		13'b1000110110101: data <= 8'b11111111;
		13'b1000110110110: data <= 8'b11111111;
		13'b1000110110111: data <= 8'b11111111;
		13'b1000110111000: data <= 8'b11111111;
		13'b1000110111001: data <= 8'b11111111;
		13'b1000111100111: data <= 8'b11111111;
		13'b1000111101000: data <= 8'b11111111;
		13'b1000111101001: data <= 8'b11111111;
		13'b1000111101010: data <= 8'b11111111;
		13'b1000111101011: data <= 8'b11111111;
		13'b1001000000100: data <= 8'b11111111;
		13'b1001000000101: data <= 8'b11111111;
		13'b1001000000110: data <= 8'b11111111;
		13'b1001000000111: data <= 8'b11111111;
		13'b1001000001000: data <= 8'b11111111;
		13'b1001000111000: data <= 8'b11111111;
		13'b1001000111001: data <= 8'b11111111;
		13'b1001000111010: data <= 8'b11111111;
		13'b1001000111011: data <= 8'b11111111;
		13'b1001000111100: data <= 8'b11111111;
		13'b1001001010011: data <= 8'b11111111;
		13'b1001001010100: data <= 8'b11111111;
		13'b1001001010101: data <= 8'b11111111;
		13'b1001001010110: data <= 8'b11111111;
		13'b1001001010111: data <= 8'b11111111;
		13'b1001010001001: data <= 8'b11111111;
		13'b1001010001010: data <= 8'b11111111;
		13'b1001010001011: data <= 8'b11111111;
		13'b1001010001100: data <= 8'b11111111;
		13'b1001010001101: data <= 8'b11111111;
		13'b1001010100010: data <= 8'b11111111;
		13'b1001010100011: data <= 8'b11111111;
		13'b1001010100100: data <= 8'b11111111;
		13'b1001010100101: data <= 8'b11111111;
		13'b1001010100110: data <= 8'b11111111;
		13'b1001011011010: data <= 8'b11111111;
		13'b1001011011011: data <= 8'b11111111;
		13'b1001011011100: data <= 8'b11111111;
		13'b1001011011101: data <= 8'b11111111;
		13'b1001011011110: data <= 8'b11111111;
		13'b1001011110001: data <= 8'b11111111;
		13'b1001011110010: data <= 8'b11111111;
		13'b1001011110011: data <= 8'b11111111;
		13'b1001011110100: data <= 8'b11111111;
		13'b1001011110101: data <= 8'b11111111;
		13'b1001100101011: data <= 8'b11111111;
		13'b1001100101100: data <= 8'b11111111;
		13'b1001100101101: data <= 8'b11111111;
		13'b1001100101110: data <= 8'b11111111;
		13'b1001100101111: data <= 8'b11111111;
		13'b1001101000000: data <= 8'b11111111;
		13'b1001101000001: data <= 8'b11111111;
		13'b1001101000010: data <= 8'b11111111;
		13'b1001101000011: data <= 8'b11111111;
		13'b1001101000100: data <= 8'b11111111;
		13'b1001101111100: data <= 8'b11111111;
		13'b1001101111101: data <= 8'b11111111;
		13'b1001101111110: data <= 8'b11111111;
		13'b1001101111111: data <= 8'b11111111;
		13'b1001110000000: data <= 8'b11111111;
		13'b1001110000001: data <= 8'b11111111;
		13'b1001110000010: data <= 8'b11111111;
		13'b1001110000011: data <= 8'b11111111;
		13'b1001110000100: data <= 8'b11111111;
		13'b1001110000101: data <= 8'b11111111;
		13'b1001110000110: data <= 8'b11111111;
		13'b1001110000111: data <= 8'b11111111;
		13'b1001110001000: data <= 8'b11111111;
		13'b1001110001001: data <= 8'b11111111;
		13'b1001110001010: data <= 8'b11111111;
		13'b1001110001011: data <= 8'b11111111;
		13'b1001110001100: data <= 8'b11111111;
		13'b1001110001101: data <= 8'b11111111;
		13'b1001110001110: data <= 8'b11111111;
		13'b1001110001111: data <= 8'b11111111;
		13'b1001110010000: data <= 8'b11111111;
		13'b1001110010001: data <= 8'b11111111;
		13'b1001110010010: data <= 8'b11111111;
		13'b1001110010011: data <= 8'b11111111;
		13'b1001111001101: data <= 8'b11111111;
		13'b1001111001110: data <= 8'b11111111;
		13'b1001111001111: data <= 8'b11111111;
		13'b1001111010000: data <= 8'b11111111;
		13'b1001111010001: data <= 8'b11111111;
		13'b1001111010010: data <= 8'b11111111;
		13'b1001111010011: data <= 8'b11111111;
		13'b1001111010100: data <= 8'b11111111;
		13'b1001111010101: data <= 8'b11111111;
		13'b1001111010110: data <= 8'b11111111;
		13'b1001111010111: data <= 8'b11111111;
		13'b1001111011000: data <= 8'b11111111;
		13'b1001111011001: data <= 8'b11111111;
		13'b1001111011010: data <= 8'b11111111;
		13'b1001111011011: data <= 8'b11111111;
		13'b1001111011100: data <= 8'b11111111;
		13'b1001111011101: data <= 8'b11111111;
		13'b1001111011110: data <= 8'b11111111;
		13'b1001111011111: data <= 8'b11111111;
		13'b1001111100000: data <= 8'b11111111;
		13'b1001111100001: data <= 8'b11111111;
		13'b1001111100010: data <= 8'b11111111;
		13'b1010000011110: data <= 8'b11111111;
		13'b1010000011111: data <= 8'b11111111;
		13'b1010000100000: data <= 8'b11111111;
		13'b1010000100001: data <= 8'b11111111;
		13'b1010000100010: data <= 8'b11111111;
		13'b1010000100011: data <= 8'b11111111;
		13'b1010000100100: data <= 8'b11111111;
		13'b1010000100101: data <= 8'b11111111;
		13'b1010000100110: data <= 8'b11111111;
		13'b1010000100111: data <= 8'b11111111;
		13'b1010000101000: data <= 8'b11111111;
		13'b1010000101001: data <= 8'b11111111;
		13'b1010000101010: data <= 8'b11111111;
		13'b1010000101011: data <= 8'b11111111;
		13'b1010000101100: data <= 8'b11111111;
		13'b1010000101101: data <= 8'b11111111;
		13'b1010000101110: data <= 8'b11111111;
		13'b1010000101111: data <= 8'b11111111;
		13'b1010000110000: data <= 8'b11111111;
		13'b1010000110001: data <= 8'b11111111;
		13'b1010001101111: data <= 8'b11111111;
		13'b1010001110000: data <= 8'b11111111;
		13'b1010001110001: data <= 8'b11111111;
		13'b1010001110010: data <= 8'b11111111;
		13'b1010001110011: data <= 8'b11111111;
		13'b1010001110100: data <= 8'b11111111;
		13'b1010001110101: data <= 8'b11111111;
		13'b1010001110110: data <= 8'b11111111;
		13'b1010001110111: data <= 8'b11111111;
		13'b1010001111000: data <= 8'b11111111;
		13'b1010001111001: data <= 8'b11111111;
		13'b1010001111010: data <= 8'b11111111;
		13'b1010001111011: data <= 8'b11111111;
		13'b1010001111100: data <= 8'b11111111;
		13'b1010001111101: data <= 8'b11111111;
		13'b1010001111110: data <= 8'b11111111;
		13'b1010001111111: data <= 8'b11111111;
		13'b1010010000000: data <= 8'b11111111;
		default: data <= 8'b00000000;
	endcase
end

endmodule
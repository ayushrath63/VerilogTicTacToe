module cursor_rom(
//inputs
clk, addr, 
//outputs
data);

(* rom_style = "block" *)

input wire clk;
input wire [12:0] addr;
output reg [7:0] data;

reg [12:0] addr_reg;

always @ (posedge clk)
	addr_reg <= addr;

always @ (*)
begin
	case(addr)
		13'b0000111100111: data <= 8'b00000011;
		13'b0000111101000: data <= 8'b00000011;
		13'b0000111101001: data <= 8'b00000011;
		13'b0000111101010: data <= 8'b00000011;
		13'b0000111101011: data <= 8'b00000011;
		13'b0000111101100: data <= 8'b00000011;
		13'b0000111101101: data <= 8'b00000011;
		13'b0000111101110: data <= 8'b00000011;
		13'b0000111101111: data <= 8'b00000011;
		13'b0000111110000: data <= 8'b00000011;
		13'b0000111110001: data <= 8'b00000011;
		13'b0000111110010: data <= 8'b00000011;
		13'b0000111110011: data <= 8'b00000011;
		13'b0000111110100: data <= 8'b00000011;
		13'b0000111110101: data <= 8'b00000011;
		13'b0000111110110: data <= 8'b00000011;
		13'b0000111110111: data <= 8'b00000011;
		13'b0000111111000: data <= 8'b00000011;
		13'b0000111111001: data <= 8'b00000011;
		13'b0000111111010: data <= 8'b00000011;
		13'b0000111111011: data <= 8'b00000011;
		13'b0000111111100: data <= 8'b00000011;
		13'b0000111111101: data <= 8'b00000011;
		13'b0000111111110: data <= 8'b00000011;
		13'b0000111111111: data <= 8'b00000011;
		13'b0001000000000: data <= 8'b00000011;
		13'b0001000001111: data <= 8'b00000011;
		13'b0001000010000: data <= 8'b00000011;
		13'b0001000010001: data <= 8'b00000011;
		13'b0001000010010: data <= 8'b00000011;
		13'b0001000010011: data <= 8'b00000011;
		13'b0001000010100: data <= 8'b00000011;
		13'b0001000010101: data <= 8'b00000011;
		13'b0001000010110: data <= 8'b00000011;
		13'b0001000010111: data <= 8'b00000011;
		13'b0001000011000: data <= 8'b00000011;
		13'b0001000011001: data <= 8'b00000011;
		13'b0001000011010: data <= 8'b00000011;
		13'b0001000011011: data <= 8'b00000011;
		13'b0001000011100: data <= 8'b00000011;
		13'b0001000011101: data <= 8'b00000011;
		13'b0001000011110: data <= 8'b00000011;
		13'b0001000011111: data <= 8'b00000011;
		13'b0001000100000: data <= 8'b00000011;
		13'b0001000100001: data <= 8'b00000011;
		13'b0001000100010: data <= 8'b00000011;
		13'b0001000100011: data <= 8'b00000011;
		13'b0001000100100: data <= 8'b00000011;
		13'b0001000100101: data <= 8'b00000011;
		13'b0001000100110: data <= 8'b00000011;
		13'b0001000100111: data <= 8'b00000011;
		13'b0001000101000: data <= 8'b00000011;
		13'b0001000110110: data <= 8'b00000011;
		13'b0001000110111: data <= 8'b00000011;
		13'b0001000111000: data <= 8'b00000011;
		13'b0001000111001: data <= 8'b00000011;
		13'b0001000111010: data <= 8'b00000011;
		13'b0001000111011: data <= 8'b00000011;
		13'b0001000111100: data <= 8'b00000011;
		13'b0001000111101: data <= 8'b00000011;
		13'b0001000111110: data <= 8'b00000011;
		13'b0001000111111: data <= 8'b00000011;
		13'b0001001000000: data <= 8'b00000011;
		13'b0001001000001: data <= 8'b00000011;
		13'b0001001000010: data <= 8'b00000011;
		13'b0001001000011: data <= 8'b00000011;
		13'b0001001000100: data <= 8'b00000011;
		13'b0001001000101: data <= 8'b00000011;
		13'b0001001000110: data <= 8'b00000011;
		13'b0001001000111: data <= 8'b00000011;
		13'b0001001001000: data <= 8'b00000011;
		13'b0001001001001: data <= 8'b00000011;
		13'b0001001001010: data <= 8'b00000011;
		13'b0001001001011: data <= 8'b00000011;
		13'b0001001001100: data <= 8'b00000011;
		13'b0001001001101: data <= 8'b00000011;
		13'b0001001001110: data <= 8'b00000011;
		13'b0001001001111: data <= 8'b00000011;
		13'b0001001010000: data <= 8'b00000011;
		13'b0001001010001: data <= 8'b00000011;
		13'b0001001011110: data <= 8'b00000011;
		13'b0001001011111: data <= 8'b00000011;
		13'b0001001100000: data <= 8'b00000011;
		13'b0001001100001: data <= 8'b00000011;
		13'b0001001100010: data <= 8'b00000011;
		13'b0001001100011: data <= 8'b00000011;
		13'b0001001100100: data <= 8'b00000011;
		13'b0001001100101: data <= 8'b00000011;
		13'b0001001100110: data <= 8'b00000011;
		13'b0001001100111: data <= 8'b00000011;
		13'b0001001101000: data <= 8'b00000011;
		13'b0001001101001: data <= 8'b00000011;
		13'b0001001101010: data <= 8'b00000011;
		13'b0001001101011: data <= 8'b00000011;
		13'b0001001101100: data <= 8'b00000011;
		13'b0001001101101: data <= 8'b00000011;
		13'b0001001101110: data <= 8'b00000011;
		13'b0001001101111: data <= 8'b00000011;
		13'b0001001110000: data <= 8'b00000011;
		13'b0001001110001: data <= 8'b00000011;
		13'b0001001110010: data <= 8'b00000011;
		13'b0001001110011: data <= 8'b00000011;
		13'b0001001110100: data <= 8'b00000011;
		13'b0001001110101: data <= 8'b00000011;
		13'b0001001110110: data <= 8'b00000011;
		13'b0001001110111: data <= 8'b00000011;
		13'b0001001111000: data <= 8'b00000011;
		13'b0001001111001: data <= 8'b00000011;
		13'b0001010000110: data <= 8'b00000011;
		13'b0001010000111: data <= 8'b00000011;
		13'b0001010001000: data <= 8'b00000011;
		13'b0001010001001: data <= 8'b00000011;
		13'b0001010001010: data <= 8'b00000011;
		13'b0001010001011: data <= 8'b00000011;
		13'b0001010001100: data <= 8'b00000011;
		13'b0001010001101: data <= 8'b00000011;
		13'b0001010001110: data <= 8'b00000011;
		13'b0001010001111: data <= 8'b00000011;
		13'b0001010010000: data <= 8'b00000011;
		13'b0001010010001: data <= 8'b00000011;
		13'b0001010010010: data <= 8'b00000011;
		13'b0001010010011: data <= 8'b00000011;
		13'b0001010010100: data <= 8'b00000011;
		13'b0001010010101: data <= 8'b00000011;
		13'b0001010010110: data <= 8'b00000011;
		13'b0001010010111: data <= 8'b00000011;
		13'b0001010011000: data <= 8'b00000011;
		13'b0001010011001: data <= 8'b00000011;
		13'b0001010011010: data <= 8'b00000011;
		13'b0001010011011: data <= 8'b00000011;
		13'b0001010011100: data <= 8'b00000011;
		13'b0001010011101: data <= 8'b00000011;
		13'b0001010011110: data <= 8'b00000011;
		13'b0001010011111: data <= 8'b00000011;
		13'b0001010100000: data <= 8'b00000011;
		13'b0001010100001: data <= 8'b00000011;
		13'b0001010101110: data <= 8'b00000011;
		13'b0001010101111: data <= 8'b00000011;
		13'b0001010110000: data <= 8'b00000011;
		13'b0001010110001: data <= 8'b00000011;
		13'b0001010110010: data <= 8'b00000011;
		13'b0001010110011: data <= 8'b00000011;
		13'b0001010110100: data <= 8'b00000011;
		13'b0001010110101: data <= 8'b00000011;
		13'b0001010110110: data <= 8'b00000011;
		13'b0001010110111: data <= 8'b00000011;
		13'b0001010111000: data <= 8'b00000011;
		13'b0001010111001: data <= 8'b00000011;
		13'b0001010111010: data <= 8'b00000011;
		13'b0001010111011: data <= 8'b00000011;
		13'b0001010111100: data <= 8'b00000011;
		13'b0001010111101: data <= 8'b00000011;
		13'b0001010111110: data <= 8'b00000011;
		13'b0001010111111: data <= 8'b00000011;
		13'b0001011000000: data <= 8'b00000011;
		13'b0001011000001: data <= 8'b00000011;
		13'b0001011000010: data <= 8'b00000011;
		13'b0001011000011: data <= 8'b00000011;
		13'b0001011000100: data <= 8'b00000011;
		13'b0001011000101: data <= 8'b00000011;
		13'b0001011000110: data <= 8'b00000011;
		13'b0001011000111: data <= 8'b00000011;
		13'b0001011001000: data <= 8'b00000011;
		13'b0001011001001: data <= 8'b00000011;
		13'b0001011010110: data <= 8'b00000011;
		13'b0001011010111: data <= 8'b00000011;
		13'b0001011011000: data <= 8'b00000011;
		13'b0001011011001: data <= 8'b00000011;
		13'b0001011011010: data <= 8'b00000011;
		13'b0001011011011: data <= 8'b00000011;
		13'b0001011011100: data <= 8'b00000011;
		13'b0001011011101: data <= 8'b00000011;
		13'b0001011011110: data <= 8'b00000011;
		13'b0001011011111: data <= 8'b00000011;
		13'b0001011100000: data <= 8'b00000011;
		13'b0001011100001: data <= 8'b00000011;
		13'b0001011100010: data <= 8'b00000011;
		13'b0001011100011: data <= 8'b00000011;
		13'b0001011100100: data <= 8'b00000011;
		13'b0001011100101: data <= 8'b00000011;
		13'b0001011100110: data <= 8'b00000011;
		13'b0001011100111: data <= 8'b00000011;
		13'b0001011101000: data <= 8'b00000011;
		13'b0001011101001: data <= 8'b00000011;
		13'b0001011101010: data <= 8'b00000011;
		13'b0001011101011: data <= 8'b00000011;
		13'b0001011101100: data <= 8'b00000011;
		13'b0001011101101: data <= 8'b00000011;
		13'b0001011101110: data <= 8'b00000011;
		13'b0001011101111: data <= 8'b00000011;
		13'b0001011110000: data <= 8'b00000011;
		13'b0001011111111: data <= 8'b00000011;
		13'b0001100000000: data <= 8'b00000011;
		13'b0001100000001: data <= 8'b00000011;
		13'b0001100000010: data <= 8'b00000011;
		13'b0001100000011: data <= 8'b00000011;
		13'b0001100000100: data <= 8'b00000011;
		13'b0001100000101: data <= 8'b00000011;
		13'b0001100000110: data <= 8'b00000011;
		13'b0001100000111: data <= 8'b00000011;
		13'b0001100001000: data <= 8'b00000011;
		13'b0001100001001: data <= 8'b00000011;
		13'b0001100001010: data <= 8'b00000011;
		13'b0001100001011: data <= 8'b00000011;
		13'b0001100001100: data <= 8'b00000011;
		13'b0001100001101: data <= 8'b00000011;
		13'b0001100001110: data <= 8'b00000011;
		13'b0001100001111: data <= 8'b00000011;
		13'b0001100010000: data <= 8'b00000011;
		13'b0001100010001: data <= 8'b00000011;
		13'b0001100010010: data <= 8'b00000011;
		13'b0001100010011: data <= 8'b00000011;
		13'b0001100010100: data <= 8'b00000011;
		13'b0001100010101: data <= 8'b00000011;
		13'b0001100010110: data <= 8'b00000011;
		13'b0001100010111: data <= 8'b00000011;
		13'b0001100011000: data <= 8'b00000011;
		13'b0001100011001: data <= 8'b00000011;
		13'b0001100100110: data <= 8'b00000011;
		13'b0001100100111: data <= 8'b00000011;
		13'b0001100101000: data <= 8'b00000011;
		13'b0001100101001: data <= 8'b00000011;
		13'b0001101100110: data <= 8'b00000011;
		13'b0001101100111: data <= 8'b00000011;
		13'b0001101101000: data <= 8'b00000011;
		13'b0001101101001: data <= 8'b00000011;
		13'b0001101110110: data <= 8'b00000011;
		13'b0001101110111: data <= 8'b00000011;
		13'b0001101111000: data <= 8'b00000011;
		13'b0001101111001: data <= 8'b00000011;
		13'b0001110110110: data <= 8'b00000011;
		13'b0001110110111: data <= 8'b00000011;
		13'b0001110111000: data <= 8'b00000011;
		13'b0001110111001: data <= 8'b00000011;
		13'b0001111000110: data <= 8'b00000011;
		13'b0001111000111: data <= 8'b00000011;
		13'b0001111001000: data <= 8'b00000011;
		13'b0001111001001: data <= 8'b00000011;
		13'b0010000000110: data <= 8'b00000011;
		13'b0010000000111: data <= 8'b00000011;
		13'b0010000001000: data <= 8'b00000011;
		13'b0010000001001: data <= 8'b00000011;
		13'b0010000010110: data <= 8'b00000011;
		13'b0010000010111: data <= 8'b00000011;
		13'b0010000011000: data <= 8'b00000011;
		13'b0010000011001: data <= 8'b00000011;
		13'b0010001010110: data <= 8'b00000011;
		13'b0010001010111: data <= 8'b00000011;
		13'b0010001011000: data <= 8'b00000011;
		13'b0010001011001: data <= 8'b00000011;
		13'b0010001100110: data <= 8'b00000011;
		13'b0010001100111: data <= 8'b00000011;
		13'b0010001101000: data <= 8'b00000011;
		13'b0010001101001: data <= 8'b00000011;
		13'b0010010100110: data <= 8'b00000011;
		13'b0010010100111: data <= 8'b00000011;
		13'b0010010101000: data <= 8'b00000011;
		13'b0010010101001: data <= 8'b00000011;
		13'b0010010110110: data <= 8'b00000011;
		13'b0010010110111: data <= 8'b00000011;
		13'b0010010111000: data <= 8'b00000011;
		13'b0010010111001: data <= 8'b00000011;
		13'b0010011110110: data <= 8'b00000011;
		13'b0010011110111: data <= 8'b00000011;
		13'b0010011111000: data <= 8'b00000011;
		13'b0010011111001: data <= 8'b00000011;
		13'b0010100000110: data <= 8'b00000011;
		13'b0010100000111: data <= 8'b00000011;
		13'b0010100001000: data <= 8'b00000011;
		13'b0010100001001: data <= 8'b00000011;
		13'b0010101000110: data <= 8'b00000011;
		13'b0010101000111: data <= 8'b00000011;
		13'b0010101001000: data <= 8'b00000011;
		13'b0010101001001: data <= 8'b00000011;
		13'b0010101010110: data <= 8'b00000011;
		13'b0010101010111: data <= 8'b00000011;
		13'b0010101011000: data <= 8'b00000011;
		13'b0010101011001: data <= 8'b00000011;
		13'b0010110010110: data <= 8'b00000011;
		13'b0010110010111: data <= 8'b00000011;
		13'b0010110011000: data <= 8'b00000011;
		13'b0010110011001: data <= 8'b00000011;
		13'b0010110100110: data <= 8'b00000011;
		13'b0010110100111: data <= 8'b00000011;
		13'b0010110101000: data <= 8'b00000011;
		13'b0010110101001: data <= 8'b00000011;
		13'b0010111100110: data <= 8'b00000011;
		13'b0010111100111: data <= 8'b00000011;
		13'b0010111101000: data <= 8'b00000011;
		13'b0010111101001: data <= 8'b00000011;
		13'b0010111110110: data <= 8'b00000011;
		13'b0010111110111: data <= 8'b00000011;
		13'b0010111111000: data <= 8'b00000011;
		13'b0010111111001: data <= 8'b00000011;
		13'b0011000110110: data <= 8'b00000011;
		13'b0011000110111: data <= 8'b00000011;
		13'b0011000111000: data <= 8'b00000011;
		13'b0011000111001: data <= 8'b00000011;
		13'b0011001000110: data <= 8'b00000011;
		13'b0011001000111: data <= 8'b00000011;
		13'b0011001001000: data <= 8'b00000011;
		13'b0011001001001: data <= 8'b00000011;
		13'b0011010000110: data <= 8'b00000011;
		13'b0011010000111: data <= 8'b00000011;
		13'b0011010001000: data <= 8'b00000011;
		13'b0011010001001: data <= 8'b00000011;
		13'b0011010010110: data <= 8'b00000011;
		13'b0011010010111: data <= 8'b00000011;
		13'b0011010011000: data <= 8'b00000011;
		13'b0011010011001: data <= 8'b00000011;
		13'b0011011010110: data <= 8'b00000011;
		13'b0011011010111: data <= 8'b00000011;
		13'b0011011011000: data <= 8'b00000011;
		13'b0011011011001: data <= 8'b00000011;
		13'b0011011100110: data <= 8'b00000011;
		13'b0011011100111: data <= 8'b00000011;
		13'b0011011101000: data <= 8'b00000011;
		13'b0011011101001: data <= 8'b00000011;
		13'b0011100100110: data <= 8'b00000011;
		13'b0011100100111: data <= 8'b00000011;
		13'b0011100101000: data <= 8'b00000011;
		13'b0011100101001: data <= 8'b00000011;
		13'b0011100110110: data <= 8'b00000011;
		13'b0011100110111: data <= 8'b00000011;
		13'b0011100111000: data <= 8'b00000011;
		13'b0011100111001: data <= 8'b00000011;
		13'b0011101110110: data <= 8'b00000011;
		13'b0011101110111: data <= 8'b00000011;
		13'b0011101111000: data <= 8'b00000011;
		13'b0011101111001: data <= 8'b00000011;
		13'b0011110000110: data <= 8'b00000011;
		13'b0011110000111: data <= 8'b00000011;
		13'b0011110001000: data <= 8'b00000011;
		13'b0011110001001: data <= 8'b00000011;
		13'b0011111000110: data <= 8'b00000011;
		13'b0011111000111: data <= 8'b00000011;
		13'b0011111001000: data <= 8'b00000011;
		13'b0011111001001: data <= 8'b00000011;
		13'b0011111010110: data <= 8'b00000011;
		13'b0011111010111: data <= 8'b00000011;
		13'b0011111011000: data <= 8'b00000011;
		13'b0011111011001: data <= 8'b00000011;
		13'b0100000010110: data <= 8'b00000011;
		13'b0100000010111: data <= 8'b00000011;
		13'b0100000011000: data <= 8'b00000011;
		13'b0100000011001: data <= 8'b00000011;
		13'b0100000100110: data <= 8'b00000011;
		13'b0100000100111: data <= 8'b00000011;
		13'b0100000101000: data <= 8'b00000011;
		13'b0100000101001: data <= 8'b00000011;
		13'b0100001100110: data <= 8'b00000011;
		13'b0100001100111: data <= 8'b00000011;
		13'b0100001101000: data <= 8'b00000011;
		13'b0100001101001: data <= 8'b00000011;
		13'b0100001110110: data <= 8'b00000011;
		13'b0100001110111: data <= 8'b00000011;
		13'b0100001111000: data <= 8'b00000011;
		13'b0100001111001: data <= 8'b00000011;
		13'b0100010110110: data <= 8'b00000011;
		13'b0100010110111: data <= 8'b00000011;
		13'b0100010111000: data <= 8'b00000011;
		13'b0100010111001: data <= 8'b00000011;
		13'b0100011000110: data <= 8'b00000011;
		13'b0100011000111: data <= 8'b00000011;
		13'b0100011001000: data <= 8'b00000011;
		13'b0100011001001: data <= 8'b00000011;
		13'b0100100000110: data <= 8'b00000011;
		13'b0100100000111: data <= 8'b00000011;
		13'b0100100001000: data <= 8'b00000011;
		13'b0100100001001: data <= 8'b00000011;
		13'b0100100010110: data <= 8'b00000011;
		13'b0100100010111: data <= 8'b00000011;
		13'b0100100011000: data <= 8'b00000011;
		13'b0100100011001: data <= 8'b00000011;
		13'b0100101010110: data <= 8'b00000011;
		13'b0100101010111: data <= 8'b00000011;
		13'b0100101011000: data <= 8'b00000011;
		13'b0100101011001: data <= 8'b00000011;
		13'b0100101100110: data <= 8'b00000011;
		13'b0100101100111: data <= 8'b00000011;
		13'b0100101101000: data <= 8'b00000011;
		13'b0100101101001: data <= 8'b00000011;
		13'b0100110100110: data <= 8'b00000011;
		13'b0100110100111: data <= 8'b00000011;
		13'b0100110101000: data <= 8'b00000011;
		13'b0100110101001: data <= 8'b00000011;
		13'b0100110110110: data <= 8'b00000011;
		13'b0100110110111: data <= 8'b00000011;
		13'b0100110111000: data <= 8'b00000011;
		13'b0100110111001: data <= 8'b00000011;
		13'b0100111110110: data <= 8'b00000011;
		13'b0100111110111: data <= 8'b00000011;
		13'b0100111111000: data <= 8'b00000011;
		13'b0100111111001: data <= 8'b00000011;
		13'b0101000000110: data <= 8'b00000011;
		13'b0101000000111: data <= 8'b00000011;
		13'b0101000001000: data <= 8'b00000011;
		13'b0101000001001: data <= 8'b00000011;
		13'b0101001000110: data <= 8'b00000011;
		13'b0101001000111: data <= 8'b00000011;
		13'b0101001001000: data <= 8'b00000011;
		13'b0101001001001: data <= 8'b00000011;
		13'b0101001010111: data <= 8'b00000011;
		13'b0101001011000: data <= 8'b00000011;
		13'b0101010010111: data <= 8'b00000011;
		13'b0101010011000: data <= 8'b00000011;
		13'b0111001100111: data <= 8'b00000011;
		13'b0111001101000: data <= 8'b00000011;
		13'b0111010100111: data <= 8'b00000011;
		13'b0111010101000: data <= 8'b00000011;
		13'b0111010110110: data <= 8'b00000011;
		13'b0111010110111: data <= 8'b00000011;
		13'b0111010111000: data <= 8'b00000011;
		13'b0111010111001: data <= 8'b00000011;
		13'b0111011110110: data <= 8'b00000011;
		13'b0111011110111: data <= 8'b00000011;
		13'b0111011111000: data <= 8'b00000011;
		13'b0111011111001: data <= 8'b00000011;
		13'b0111100000110: data <= 8'b00000011;
		13'b0111100000111: data <= 8'b00000011;
		13'b0111100001000: data <= 8'b00000011;
		13'b0111100001001: data <= 8'b00000011;
		13'b0111101000110: data <= 8'b00000011;
		13'b0111101000111: data <= 8'b00000011;
		13'b0111101001000: data <= 8'b00000011;
		13'b0111101001001: data <= 8'b00000011;
		13'b0111101010110: data <= 8'b00000011;
		13'b0111101010111: data <= 8'b00000011;
		13'b0111101011000: data <= 8'b00000011;
		13'b0111101011001: data <= 8'b00000011;
		13'b0111110010110: data <= 8'b00000011;
		13'b0111110010111: data <= 8'b00000011;
		13'b0111110011000: data <= 8'b00000011;
		13'b0111110011001: data <= 8'b00000011;
		13'b0111110100110: data <= 8'b00000011;
		13'b0111110100111: data <= 8'b00000011;
		13'b0111110101000: data <= 8'b00000011;
		13'b0111110101001: data <= 8'b00000011;
		13'b0111111100110: data <= 8'b00000011;
		13'b0111111100111: data <= 8'b00000011;
		13'b0111111101000: data <= 8'b00000011;
		13'b0111111101001: data <= 8'b00000011;
		13'b0111111110110: data <= 8'b00000011;
		13'b0111111110111: data <= 8'b00000011;
		13'b0111111111000: data <= 8'b00000011;
		13'b0111111111001: data <= 8'b00000011;
		13'b1000000110110: data <= 8'b00000011;
		13'b1000000110111: data <= 8'b00000011;
		13'b1000000111000: data <= 8'b00000011;
		13'b1000000111001: data <= 8'b00000011;
		13'b1000001000110: data <= 8'b00000011;
		13'b1000001000111: data <= 8'b00000011;
		13'b1000001001000: data <= 8'b00000011;
		13'b1000001001001: data <= 8'b00000011;
		13'b1000010000110: data <= 8'b00000011;
		13'b1000010000111: data <= 8'b00000011;
		13'b1000010001000: data <= 8'b00000011;
		13'b1000010001001: data <= 8'b00000011;
		13'b1000010010110: data <= 8'b00000011;
		13'b1000010010111: data <= 8'b00000011;
		13'b1000010011000: data <= 8'b00000011;
		13'b1000010011001: data <= 8'b00000011;
		13'b1000011010110: data <= 8'b00000011;
		13'b1000011010111: data <= 8'b00000011;
		13'b1000011011000: data <= 8'b00000011;
		13'b1000011011001: data <= 8'b00000011;
		13'b1000011100110: data <= 8'b00000011;
		13'b1000011100111: data <= 8'b00000011;
		13'b1000011101000: data <= 8'b00000011;
		13'b1000011101001: data <= 8'b00000011;
		13'b1000100100110: data <= 8'b00000011;
		13'b1000100100111: data <= 8'b00000011;
		13'b1000100101000: data <= 8'b00000011;
		13'b1000100101001: data <= 8'b00000011;
		13'b1000100110110: data <= 8'b00000011;
		13'b1000100110111: data <= 8'b00000011;
		13'b1000100111000: data <= 8'b00000011;
		13'b1000100111001: data <= 8'b00000011;
		13'b1000101110110: data <= 8'b00000011;
		13'b1000101110111: data <= 8'b00000011;
		13'b1000101111000: data <= 8'b00000011;
		13'b1000101111001: data <= 8'b00000011;
		13'b1000110000110: data <= 8'b00000011;
		13'b1000110000111: data <= 8'b00000011;
		13'b1000110001000: data <= 8'b00000011;
		13'b1000110001001: data <= 8'b00000011;
		13'b1000111000110: data <= 8'b00000011;
		13'b1000111000111: data <= 8'b00000011;
		13'b1000111001000: data <= 8'b00000011;
		13'b1000111001001: data <= 8'b00000011;
		13'b1000111010110: data <= 8'b00000011;
		13'b1000111010111: data <= 8'b00000011;
		13'b1000111011000: data <= 8'b00000011;
		13'b1000111011001: data <= 8'b00000011;
		13'b1001000010110: data <= 8'b00000011;
		13'b1001000010111: data <= 8'b00000011;
		13'b1001000011000: data <= 8'b00000011;
		13'b1001000011001: data <= 8'b00000011;
		13'b1001000100110: data <= 8'b00000011;
		13'b1001000100111: data <= 8'b00000011;
		13'b1001000101000: data <= 8'b00000011;
		13'b1001000101001: data <= 8'b00000011;
		13'b1001001100110: data <= 8'b00000011;
		13'b1001001100111: data <= 8'b00000011;
		13'b1001001101000: data <= 8'b00000011;
		13'b1001001101001: data <= 8'b00000011;
		13'b1001001110110: data <= 8'b00000011;
		13'b1001001110111: data <= 8'b00000011;
		13'b1001001111000: data <= 8'b00000011;
		13'b1001001111001: data <= 8'b00000011;
		13'b1001010110110: data <= 8'b00000011;
		13'b1001010110111: data <= 8'b00000011;
		13'b1001010111000: data <= 8'b00000011;
		13'b1001010111001: data <= 8'b00000011;
		13'b1001011000110: data <= 8'b00000011;
		13'b1001011000111: data <= 8'b00000011;
		13'b1001011001000: data <= 8'b00000011;
		13'b1001011001001: data <= 8'b00000011;
		13'b1001100000110: data <= 8'b00000011;
		13'b1001100000111: data <= 8'b00000011;
		13'b1001100001000: data <= 8'b00000011;
		13'b1001100001001: data <= 8'b00000011;
		13'b1001100010110: data <= 8'b00000011;
		13'b1001100010111: data <= 8'b00000011;
		13'b1001100011000: data <= 8'b00000011;
		13'b1001100011001: data <= 8'b00000011;
		13'b1001101010110: data <= 8'b00000011;
		13'b1001101010111: data <= 8'b00000011;
		13'b1001101011000: data <= 8'b00000011;
		13'b1001101011001: data <= 8'b00000011;
		13'b1001101100110: data <= 8'b00000011;
		13'b1001101100111: data <= 8'b00000011;
		13'b1001101101000: data <= 8'b00000011;
		13'b1001101101001: data <= 8'b00000011;
		13'b1001110100110: data <= 8'b00000011;
		13'b1001110100111: data <= 8'b00000011;
		13'b1001110101000: data <= 8'b00000011;
		13'b1001110101001: data <= 8'b00000011;
		13'b1001110110110: data <= 8'b00000011;
		13'b1001110110111: data <= 8'b00000011;
		13'b1001110111000: data <= 8'b00000011;
		13'b1001110111001: data <= 8'b00000011;
		13'b1001111110110: data <= 8'b00000011;
		13'b1001111110111: data <= 8'b00000011;
		13'b1001111111000: data <= 8'b00000011;
		13'b1001111111001: data <= 8'b00000011;
		13'b1010000000110: data <= 8'b00000011;
		13'b1010000000111: data <= 8'b00000011;
		13'b1010000001000: data <= 8'b00000011;
		13'b1010000001001: data <= 8'b00000011;
		13'b1010001000110: data <= 8'b00000011;
		13'b1010001000111: data <= 8'b00000011;
		13'b1010001001000: data <= 8'b00000011;
		13'b1010001001001: data <= 8'b00000011;
		13'b1010001010110: data <= 8'b00000011;
		13'b1010001010111: data <= 8'b00000011;
		13'b1010001011000: data <= 8'b00000011;
		13'b1010001011001: data <= 8'b00000011;
		13'b1010010010110: data <= 8'b00000011;
		13'b1010010010111: data <= 8'b00000011;
		13'b1010010011000: data <= 8'b00000011;
		13'b1010010011001: data <= 8'b00000011;
		13'b1010010100110: data <= 8'b00000011;
		13'b1010010100111: data <= 8'b00000011;
		13'b1010010101000: data <= 8'b00000011;
		13'b1010010101001: data <= 8'b00000011;
		13'b1010011100110: data <= 8'b00000011;
		13'b1010011100111: data <= 8'b00000011;
		13'b1010011101000: data <= 8'b00000011;
		13'b1010011101001: data <= 8'b00000011;
		13'b1010011110110: data <= 8'b00000011;
		13'b1010011110111: data <= 8'b00000011;
		13'b1010011111000: data <= 8'b00000011;
		13'b1010011111001: data <= 8'b00000011;
		13'b1010100110110: data <= 8'b00000011;
		13'b1010100110111: data <= 8'b00000011;
		13'b1010100111000: data <= 8'b00000011;
		13'b1010100111001: data <= 8'b00000011;
		13'b1010101000110: data <= 8'b00000011;
		13'b1010101000111: data <= 8'b00000011;
		13'b1010101001000: data <= 8'b00000011;
		13'b1010101001001: data <= 8'b00000011;
		13'b1010110000110: data <= 8'b00000011;
		13'b1010110000111: data <= 8'b00000011;
		13'b1010110001000: data <= 8'b00000011;
		13'b1010110001001: data <= 8'b00000011;
		13'b1010110010110: data <= 8'b00000011;
		13'b1010110010111: data <= 8'b00000011;
		13'b1010110011000: data <= 8'b00000011;
		13'b1010110011001: data <= 8'b00000011;
		13'b1010111010110: data <= 8'b00000011;
		13'b1010111010111: data <= 8'b00000011;
		13'b1010111011000: data <= 8'b00000011;
		13'b1010111011001: data <= 8'b00000011;
		13'b1010111100110: data <= 8'b00000011;
		13'b1010111100111: data <= 8'b00000011;
		13'b1010111101000: data <= 8'b00000011;
		13'b1010111101001: data <= 8'b00000011;
		13'b1010111101010: data <= 8'b00000011;
		13'b1010111101011: data <= 8'b00000011;
		13'b1010111101100: data <= 8'b00000011;
		13'b1010111101101: data <= 8'b00000011;
		13'b1010111101110: data <= 8'b00000011;
		13'b1010111101111: data <= 8'b00000011;
		13'b1010111110000: data <= 8'b00000011;
		13'b1010111110001: data <= 8'b00000011;
		13'b1010111110010: data <= 8'b00000011;
		13'b1010111110011: data <= 8'b00000011;
		13'b1010111110100: data <= 8'b00000011;
		13'b1010111110101: data <= 8'b00000011;
		13'b1010111110110: data <= 8'b00000011;
		13'b1010111110111: data <= 8'b00000011;
		13'b1010111111000: data <= 8'b00000011;
		13'b1010111111001: data <= 8'b00000011;
		13'b1010111111010: data <= 8'b00000011;
		13'b1010111111011: data <= 8'b00000011;
		13'b1010111111100: data <= 8'b00000011;
		13'b1010111111101: data <= 8'b00000011;
		13'b1010111111110: data <= 8'b00000011;
		13'b1010111111111: data <= 8'b00000011;
		13'b1011000000000: data <= 8'b00000011;
		13'b1011000001111: data <= 8'b00000011;
		13'b1011000010000: data <= 8'b00000011;
		13'b1011000010001: data <= 8'b00000011;
		13'b1011000010010: data <= 8'b00000011;
		13'b1011000010011: data <= 8'b00000011;
		13'b1011000010100: data <= 8'b00000011;
		13'b1011000010101: data <= 8'b00000011;
		13'b1011000010110: data <= 8'b00000011;
		13'b1011000010111: data <= 8'b00000011;
		13'b1011000011000: data <= 8'b00000011;
		13'b1011000011001: data <= 8'b00000011;
		13'b1011000011010: data <= 8'b00000011;
		13'b1011000011011: data <= 8'b00000011;
		13'b1011000011100: data <= 8'b00000011;
		13'b1011000011101: data <= 8'b00000011;
		13'b1011000011110: data <= 8'b00000011;
		13'b1011000011111: data <= 8'b00000011;
		13'b1011000100000: data <= 8'b00000011;
		13'b1011000100001: data <= 8'b00000011;
		13'b1011000100010: data <= 8'b00000011;
		13'b1011000100011: data <= 8'b00000011;
		13'b1011000100100: data <= 8'b00000011;
		13'b1011000100101: data <= 8'b00000011;
		13'b1011000100110: data <= 8'b00000011;
		13'b1011000100111: data <= 8'b00000011;
		13'b1011000101000: data <= 8'b00000011;
		13'b1011000101001: data <= 8'b00000011;
		13'b1011000110110: data <= 8'b00000011;
		13'b1011000110111: data <= 8'b00000011;
		13'b1011000111000: data <= 8'b00000011;
		13'b1011000111001: data <= 8'b00000011;
		13'b1011000111010: data <= 8'b00000011;
		13'b1011000111011: data <= 8'b00000011;
		13'b1011000111100: data <= 8'b00000011;
		13'b1011000111101: data <= 8'b00000011;
		13'b1011000111110: data <= 8'b00000011;
		13'b1011000111111: data <= 8'b00000011;
		13'b1011001000000: data <= 8'b00000011;
		13'b1011001000001: data <= 8'b00000011;
		13'b1011001000010: data <= 8'b00000011;
		13'b1011001000011: data <= 8'b00000011;
		13'b1011001000100: data <= 8'b00000011;
		13'b1011001000101: data <= 8'b00000011;
		13'b1011001000110: data <= 8'b00000011;
		13'b1011001000111: data <= 8'b00000011;
		13'b1011001001000: data <= 8'b00000011;
		13'b1011001001001: data <= 8'b00000011;
		13'b1011001001010: data <= 8'b00000011;
		13'b1011001001011: data <= 8'b00000011;
		13'b1011001001100: data <= 8'b00000011;
		13'b1011001001101: data <= 8'b00000011;
		13'b1011001001110: data <= 8'b00000011;
		13'b1011001001111: data <= 8'b00000011;
		13'b1011001010000: data <= 8'b00000011;
		13'b1011001010001: data <= 8'b00000011;
		13'b1011001011110: data <= 8'b00000011;
		13'b1011001011111: data <= 8'b00000011;
		13'b1011001100000: data <= 8'b00000011;
		13'b1011001100001: data <= 8'b00000011;
		13'b1011001100010: data <= 8'b00000011;
		13'b1011001100011: data <= 8'b00000011;
		13'b1011001100100: data <= 8'b00000011;
		13'b1011001100101: data <= 8'b00000011;
		13'b1011001100110: data <= 8'b00000011;
		13'b1011001100111: data <= 8'b00000011;
		13'b1011001101000: data <= 8'b00000011;
		13'b1011001101001: data <= 8'b00000011;
		13'b1011001101010: data <= 8'b00000011;
		13'b1011001101011: data <= 8'b00000011;
		13'b1011001101100: data <= 8'b00000011;
		13'b1011001101101: data <= 8'b00000011;
		13'b1011001101110: data <= 8'b00000011;
		13'b1011001101111: data <= 8'b00000011;
		13'b1011001110000: data <= 8'b00000011;
		13'b1011001110001: data <= 8'b00000011;
		13'b1011001110010: data <= 8'b00000011;
		13'b1011001110011: data <= 8'b00000011;
		13'b1011001110100: data <= 8'b00000011;
		13'b1011001110101: data <= 8'b00000011;
		13'b1011001110110: data <= 8'b00000011;
		13'b1011001110111: data <= 8'b00000011;
		13'b1011001111000: data <= 8'b00000011;
		13'b1011001111001: data <= 8'b00000011;
		13'b1011010000110: data <= 8'b00000011;
		13'b1011010000111: data <= 8'b00000011;
		13'b1011010001000: data <= 8'b00000011;
		13'b1011010001001: data <= 8'b00000011;
		13'b1011010001010: data <= 8'b00000011;
		13'b1011010001011: data <= 8'b00000011;
		13'b1011010001100: data <= 8'b00000011;
		13'b1011010001101: data <= 8'b00000011;
		13'b1011010001110: data <= 8'b00000011;
		13'b1011010001111: data <= 8'b00000011;
		13'b1011010010000: data <= 8'b00000011;
		13'b1011010010001: data <= 8'b00000011;
		13'b1011010010010: data <= 8'b00000011;
		13'b1011010010011: data <= 8'b00000011;
		13'b1011010010100: data <= 8'b00000011;
		13'b1011010010101: data <= 8'b00000011;
		13'b1011010010110: data <= 8'b00000011;
		13'b1011010010111: data <= 8'b00000011;
		13'b1011010011000: data <= 8'b00000011;
		13'b1011010011001: data <= 8'b00000011;
		13'b1011010011010: data <= 8'b00000011;
		13'b1011010011011: data <= 8'b00000011;
		13'b1011010011100: data <= 8'b00000011;
		13'b1011010011101: data <= 8'b00000011;
		13'b1011010011110: data <= 8'b00000011;
		13'b1011010011111: data <= 8'b00000011;
		13'b1011010100000: data <= 8'b00000011;
		13'b1011010100001: data <= 8'b00000011;
		13'b1011010101110: data <= 8'b00000011;
		13'b1011010101111: data <= 8'b00000011;
		13'b1011010110000: data <= 8'b00000011;
		13'b1011010110001: data <= 8'b00000011;
		13'b1011010110010: data <= 8'b00000011;
		13'b1011010110011: data <= 8'b00000011;
		13'b1011010110100: data <= 8'b00000011;
		13'b1011010110101: data <= 8'b00000011;
		13'b1011010110110: data <= 8'b00000011;
		13'b1011010110111: data <= 8'b00000011;
		13'b1011010111000: data <= 8'b00000011;
		13'b1011010111001: data <= 8'b00000011;
		13'b1011010111010: data <= 8'b00000011;
		13'b1011010111011: data <= 8'b00000011;
		13'b1011010111100: data <= 8'b00000011;
		13'b1011010111101: data <= 8'b00000011;
		13'b1011010111110: data <= 8'b00000011;
		13'b1011010111111: data <= 8'b00000011;
		13'b1011011000000: data <= 8'b00000011;
		13'b1011011000001: data <= 8'b00000011;
		13'b1011011000010: data <= 8'b00000011;
		13'b1011011000011: data <= 8'b00000011;
		13'b1011011000100: data <= 8'b00000011;
		13'b1011011000101: data <= 8'b00000011;
		13'b1011011000110: data <= 8'b00000011;
		13'b1011011000111: data <= 8'b00000011;
		13'b1011011001000: data <= 8'b00000011;
		13'b1011011001001: data <= 8'b00000011;
		13'b1011011010111: data <= 8'b00000011;
		13'b1011011011000: data <= 8'b00000011;
		13'b1011011011001: data <= 8'b00000011;
		13'b1011011011010: data <= 8'b00000011;
		13'b1011011011011: data <= 8'b00000011;
		13'b1011011011100: data <= 8'b00000011;
		13'b1011011011101: data <= 8'b00000011;
		13'b1011011011110: data <= 8'b00000011;
		13'b1011011011111: data <= 8'b00000011;
		13'b1011011100000: data <= 8'b00000011;
		13'b1011011100001: data <= 8'b00000011;
		13'b1011011100010: data <= 8'b00000011;
		13'b1011011100011: data <= 8'b00000011;
		13'b1011011100100: data <= 8'b00000011;
		13'b1011011100101: data <= 8'b00000011;
		13'b1011011100110: data <= 8'b00000011;
		13'b1011011100111: data <= 8'b00000011;
		13'b1011011101000: data <= 8'b00000011;
		13'b1011011101001: data <= 8'b00000011;
		13'b1011011101010: data <= 8'b00000011;
		13'b1011011101011: data <= 8'b00000011;
		13'b1011011101100: data <= 8'b00000011;
		13'b1011011101101: data <= 8'b00000011;
		13'b1011011101110: data <= 8'b00000011;
		13'b1011011101111: data <= 8'b00000011;
		13'b1011011110000: data <= 8'b00000011;
		13'b1011011111111: data <= 8'b00000011;
		13'b1011100000000: data <= 8'b00000011;
		13'b1011100000001: data <= 8'b00000011;
		13'b1011100000010: data <= 8'b00000011;
		13'b1011100000011: data <= 8'b00000011;
		13'b1011100000100: data <= 8'b00000011;
		13'b1011100000101: data <= 8'b00000011;
		13'b1011100000110: data <= 8'b00000011;
		13'b1011100000111: data <= 8'b00000011;
		13'b1011100001000: data <= 8'b00000011;
		13'b1011100001001: data <= 8'b00000011;
		13'b1011100001010: data <= 8'b00000011;
		13'b1011100001011: data <= 8'b00000011;
		13'b1011100001100: data <= 8'b00000011;
		13'b1011100001101: data <= 8'b00000011;
		13'b1011100001110: data <= 8'b00000011;
		13'b1011100001111: data <= 8'b00000011;
		13'b1011100010000: data <= 8'b00000011;
		13'b1011100010001: data <= 8'b00000011;
		13'b1011100010010: data <= 8'b00000011;
		13'b1011100010011: data <= 8'b00000011;
		13'b1011100010100: data <= 8'b00000011;
		13'b1011100010101: data <= 8'b00000011;
		13'b1011100010110: data <= 8'b00000011;
		13'b1011100010111: data <= 8'b00000011;
		13'b1011100011000: data <= 8'b00000011;
		default: data <= 8'b00000000;
	endcase
end

endmodule
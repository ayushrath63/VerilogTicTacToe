module x_rom(
//inputs
clk, addr, 
//outputs
data);

(* rom_style = "block" *)

input wire clk;
input wire [12:0] addr;
output reg [7:0] data;

reg [12:0] addr_reg;

always @ (posedge clk)
	addr_reg <= addr;

always @ (*)
begin
	case(addr)
		13'b0010001101111: data <= 8'b11111111;
		13'b0010001110000: data <= 8'b11111111;
		13'b0010010011111: data <= 8'b11111111;
		13'b0010010100000: data <= 8'b11111111;
		13'b0010010111110: data <= 8'b11111111;
		13'b0010010111111: data <= 8'b11111111;
		13'b0010011000000: data <= 8'b11111111;
		13'b0010011000001: data <= 8'b11111111;
		13'b0010011101110: data <= 8'b11111111;
		13'b0010011101111: data <= 8'b11111111;
		13'b0010011110000: data <= 8'b11111111;
		13'b0010011110001: data <= 8'b11111111;
		13'b0010100001110: data <= 8'b11111111;
		13'b0010100001111: data <= 8'b11111111;
		13'b0010100010000: data <= 8'b11111111;
		13'b0010100010001: data <= 8'b11111111;
		13'b0010100010010: data <= 8'b11111111;
		13'b0010100111101: data <= 8'b11111111;
		13'b0010100111110: data <= 8'b11111111;
		13'b0010100111111: data <= 8'b11111111;
		13'b0010101000000: data <= 8'b11111111;
		13'b0010101000001: data <= 8'b11111111;
		13'b0010101011111: data <= 8'b11111111;
		13'b0010101100000: data <= 8'b11111111;
		13'b0010101100001: data <= 8'b11111111;
		13'b0010101100010: data <= 8'b11111111;
		13'b0010101100011: data <= 8'b11111111;
		13'b0010110001100: data <= 8'b11111111;
		13'b0010110001101: data <= 8'b11111111;
		13'b0010110001110: data <= 8'b11111111;
		13'b0010110001111: data <= 8'b11111111;
		13'b0010110010000: data <= 8'b11111111;
		13'b0010110110000: data <= 8'b11111111;
		13'b0010110110001: data <= 8'b11111111;
		13'b0010110110010: data <= 8'b11111111;
		13'b0010110110011: data <= 8'b11111111;
		13'b0010110110100: data <= 8'b11111111;
		13'b0010111011011: data <= 8'b11111111;
		13'b0010111011100: data <= 8'b11111111;
		13'b0010111011101: data <= 8'b11111111;
		13'b0010111011110: data <= 8'b11111111;
		13'b0010111011111: data <= 8'b11111111;
		13'b0011000000001: data <= 8'b11111111;
		13'b0011000000010: data <= 8'b11111111;
		13'b0011000000011: data <= 8'b11111111;
		13'b0011000000100: data <= 8'b11111111;
		13'b0011000000101: data <= 8'b11111111;
		13'b0011000101010: data <= 8'b11111111;
		13'b0011000101011: data <= 8'b11111111;
		13'b0011000101100: data <= 8'b11111111;
		13'b0011000101101: data <= 8'b11111111;
		13'b0011000101110: data <= 8'b11111111;
		13'b0011001010010: data <= 8'b11111111;
		13'b0011001010011: data <= 8'b11111111;
		13'b0011001010100: data <= 8'b11111111;
		13'b0011001010101: data <= 8'b11111111;
		13'b0011001010110: data <= 8'b11111111;
		13'b0011001111001: data <= 8'b11111111;
		13'b0011001111010: data <= 8'b11111111;
		13'b0011001111011: data <= 8'b11111111;
		13'b0011001111100: data <= 8'b11111111;
		13'b0011001111101: data <= 8'b11111111;
		13'b0011010100011: data <= 8'b11111111;
		13'b0011010100100: data <= 8'b11111111;
		13'b0011010100101: data <= 8'b11111111;
		13'b0011010100110: data <= 8'b11111111;
		13'b0011010100111: data <= 8'b11111111;
		13'b0011011001000: data <= 8'b11111111;
		13'b0011011001001: data <= 8'b11111111;
		13'b0011011001010: data <= 8'b11111111;
		13'b0011011001011: data <= 8'b11111111;
		13'b0011011001100: data <= 8'b11111111;
		13'b0011011110100: data <= 8'b11111111;
		13'b0011011110101: data <= 8'b11111111;
		13'b0011011110110: data <= 8'b11111111;
		13'b0011011110111: data <= 8'b11111111;
		13'b0011011111000: data <= 8'b11111111;
		13'b0011100010111: data <= 8'b11111111;
		13'b0011100011000: data <= 8'b11111111;
		13'b0011100011001: data <= 8'b11111111;
		13'b0011100011010: data <= 8'b11111111;
		13'b0011100011011: data <= 8'b11111111;
		13'b0011101000101: data <= 8'b11111111;
		13'b0011101000110: data <= 8'b11111111;
		13'b0011101000111: data <= 8'b11111111;
		13'b0011101001000: data <= 8'b11111111;
		13'b0011101001001: data <= 8'b11111111;
		13'b0011101100110: data <= 8'b11111111;
		13'b0011101100111: data <= 8'b11111111;
		13'b0011101101000: data <= 8'b11111111;
		13'b0011101101001: data <= 8'b11111111;
		13'b0011101101010: data <= 8'b11111111;
		13'b0011110010110: data <= 8'b11111111;
		13'b0011110010111: data <= 8'b11111111;
		13'b0011110011000: data <= 8'b11111111;
		13'b0011110011001: data <= 8'b11111111;
		13'b0011110011010: data <= 8'b11111111;
		13'b0011110110101: data <= 8'b11111111;
		13'b0011110110110: data <= 8'b11111111;
		13'b0011110110111: data <= 8'b11111111;
		13'b0011110111000: data <= 8'b11111111;
		13'b0011110111001: data <= 8'b11111111;
		13'b0011111100111: data <= 8'b11111111;
		13'b0011111101000: data <= 8'b11111111;
		13'b0011111101001: data <= 8'b11111111;
		13'b0011111101010: data <= 8'b11111111;
		13'b0011111101011: data <= 8'b11111111;
		13'b0100000000100: data <= 8'b11111111;
		13'b0100000000101: data <= 8'b11111111;
		13'b0100000000110: data <= 8'b11111111;
		13'b0100000000111: data <= 8'b11111111;
		13'b0100000001000: data <= 8'b11111111;
		13'b0100000111000: data <= 8'b11111111;
		13'b0100000111001: data <= 8'b11111111;
		13'b0100000111010: data <= 8'b11111111;
		13'b0100000111011: data <= 8'b11111111;
		13'b0100000111100: data <= 8'b11111111;
		13'b0100001010011: data <= 8'b11111111;
		13'b0100001010100: data <= 8'b11111111;
		13'b0100001010101: data <= 8'b11111111;
		13'b0100001010110: data <= 8'b11111111;
		13'b0100001010111: data <= 8'b11111111;
		13'b0100010001001: data <= 8'b11111111;
		13'b0100010001010: data <= 8'b11111111;
		13'b0100010001011: data <= 8'b11111111;
		13'b0100010001100: data <= 8'b11111111;
		13'b0100010001101: data <= 8'b11111111;
		13'b0100010100010: data <= 8'b11111111;
		13'b0100010100011: data <= 8'b11111111;
		13'b0100010100100: data <= 8'b11111111;
		13'b0100010100101: data <= 8'b11111111;
		13'b0100010100110: data <= 8'b11111111;
		13'b0100011011010: data <= 8'b11111111;
		13'b0100011011011: data <= 8'b11111111;
		13'b0100011011100: data <= 8'b11111111;
		13'b0100011011101: data <= 8'b11111111;
		13'b0100011011110: data <= 8'b11111111;
		13'b0100011110001: data <= 8'b11111111;
		13'b0100011110010: data <= 8'b11111111;
		13'b0100011110011: data <= 8'b11111111;
		13'b0100011110100: data <= 8'b11111111;
		13'b0100011110101: data <= 8'b11111111;
		13'b0100100101011: data <= 8'b11111111;
		13'b0100100101100: data <= 8'b11111111;
		13'b0100100101101: data <= 8'b11111111;
		13'b0100100101110: data <= 8'b11111111;
		13'b0100100101111: data <= 8'b11111111;
		13'b0100101000000: data <= 8'b11111111;
		13'b0100101000001: data <= 8'b11111111;
		13'b0100101000010: data <= 8'b11111111;
		13'b0100101000011: data <= 8'b11111111;
		13'b0100101000100: data <= 8'b11111111;
		13'b0100101111100: data <= 8'b11111111;
		13'b0100101111101: data <= 8'b11111111;
		13'b0100101111110: data <= 8'b11111111;
		13'b0100101111111: data <= 8'b11111111;
		13'b0100110000000: data <= 8'b11111111;
		13'b0100110001111: data <= 8'b11111111;
		13'b0100110010000: data <= 8'b11111111;
		13'b0100110010001: data <= 8'b11111111;
		13'b0100110010010: data <= 8'b11111111;
		13'b0100110010011: data <= 8'b11111111;
		13'b0100111001101: data <= 8'b11111111;
		13'b0100111001110: data <= 8'b11111111;
		13'b0100111001111: data <= 8'b11111111;
		13'b0100111010000: data <= 8'b11111111;
		13'b0100111010001: data <= 8'b11111111;
		13'b0100111011110: data <= 8'b11111111;
		13'b0100111011111: data <= 8'b11111111;
		13'b0100111100000: data <= 8'b11111111;
		13'b0100111100001: data <= 8'b11111111;
		13'b0100111100010: data <= 8'b11111111;
		13'b0101000011110: data <= 8'b11111111;
		13'b0101000011111: data <= 8'b11111111;
		13'b0101000100000: data <= 8'b11111111;
		13'b0101000100001: data <= 8'b11111111;
		13'b0101000100010: data <= 8'b11111111;
		13'b0101000101101: data <= 8'b11111111;
		13'b0101000101110: data <= 8'b11111111;
		13'b0101000101111: data <= 8'b11111111;
		13'b0101000110000: data <= 8'b11111111;
		13'b0101000110001: data <= 8'b11111111;
		13'b0101001101111: data <= 8'b11111111;
		13'b0101001110000: data <= 8'b11111111;
		13'b0101001110001: data <= 8'b11111111;
		13'b0101001110010: data <= 8'b11111111;
		13'b0101001110011: data <= 8'b11111111;
		13'b0101001111100: data <= 8'b11111111;
		13'b0101001111101: data <= 8'b11111111;
		13'b0101001111110: data <= 8'b11111111;
		13'b0101001111111: data <= 8'b11111111;
		13'b0101010000000: data <= 8'b11111111;
		13'b0101011000000: data <= 8'b11111111;
		13'b0101011000001: data <= 8'b11111111;
		13'b0101011000010: data <= 8'b11111111;
		13'b0101011000011: data <= 8'b11111111;
		13'b0101011000100: data <= 8'b11111111;
		13'b0101011001011: data <= 8'b11111111;
		13'b0101011001100: data <= 8'b11111111;
		13'b0101011001101: data <= 8'b11111111;
		13'b0101011001110: data <= 8'b11111111;
		13'b0101011001111: data <= 8'b11111111;
		13'b0101100010001: data <= 8'b11111111;
		13'b0101100010010: data <= 8'b11111111;
		13'b0101100010011: data <= 8'b11111111;
		13'b0101100010100: data <= 8'b11111111;
		13'b0101100010101: data <= 8'b11111111;
		13'b0101100011010: data <= 8'b11111111;
		13'b0101100011011: data <= 8'b11111111;
		13'b0101100011100: data <= 8'b11111111;
		13'b0101100011101: data <= 8'b11111111;
		13'b0101100011110: data <= 8'b11111111;
		13'b0101101100010: data <= 8'b11111111;
		13'b0101101100011: data <= 8'b11111111;
		13'b0101101100100: data <= 8'b11111111;
		13'b0101101100101: data <= 8'b11111111;
		13'b0101101100110: data <= 8'b11111111;
		13'b0101101101001: data <= 8'b11111111;
		13'b0101101101010: data <= 8'b11111111;
		13'b0101101101011: data <= 8'b11111111;
		13'b0101101101100: data <= 8'b11111111;
		13'b0101101101101: data <= 8'b11111111;
		13'b0101110110011: data <= 8'b11111111;
		13'b0101110110100: data <= 8'b11111111;
		13'b0101110110101: data <= 8'b11111111;
		13'b0101110110110: data <= 8'b11111111;
		13'b0101110110111: data <= 8'b11111111;
		13'b0101110111000: data <= 8'b11111111;
		13'b0101110111001: data <= 8'b11111111;
		13'b0101110111010: data <= 8'b11111111;
		13'b0101110111011: data <= 8'b11111111;
		13'b0101110111100: data <= 8'b11111111;
		13'b0110000000100: data <= 8'b11111111;
		13'b0110000000101: data <= 8'b11111111;
		13'b0110000000110: data <= 8'b11111111;
		13'b0110000000111: data <= 8'b11111111;
		13'b0110000001000: data <= 8'b11111111;
		13'b0110000001001: data <= 8'b11111111;
		13'b0110000001010: data <= 8'b11111111;
		13'b0110000001011: data <= 8'b11111111;
		13'b0110001010101: data <= 8'b11111111;
		13'b0110001010110: data <= 8'b11111111;
		13'b0110001010111: data <= 8'b11111111;
		13'b0110001011000: data <= 8'b11111111;
		13'b0110001011001: data <= 8'b11111111;
		13'b0110001011010: data <= 8'b11111111;
		13'b0110010100101: data <= 8'b11111111;
		13'b0110010100110: data <= 8'b11111111;
		13'b0110010100111: data <= 8'b11111111;
		13'b0110010101000: data <= 8'b11111111;
		13'b0110010101001: data <= 8'b11111111;
		13'b0110010101010: data <= 8'b11111111;
		13'b0110011110100: data <= 8'b11111111;
		13'b0110011110101: data <= 8'b11111111;
		13'b0110011110110: data <= 8'b11111111;
		13'b0110011110111: data <= 8'b11111111;
		13'b0110011111000: data <= 8'b11111111;
		13'b0110011111001: data <= 8'b11111111;
		13'b0110011111010: data <= 8'b11111111;
		13'b0110011111011: data <= 8'b11111111;
		13'b0110101000011: data <= 8'b11111111;
		13'b0110101000100: data <= 8'b11111111;
		13'b0110101000101: data <= 8'b11111111;
		13'b0110101000110: data <= 8'b11111111;
		13'b0110101000111: data <= 8'b11111111;
		13'b0110101001000: data <= 8'b11111111;
		13'b0110101001001: data <= 8'b11111111;
		13'b0110101001010: data <= 8'b11111111;
		13'b0110101001011: data <= 8'b11111111;
		13'b0110101001100: data <= 8'b11111111;
		13'b0110110010010: data <= 8'b11111111;
		13'b0110110010011: data <= 8'b11111111;
		13'b0110110010100: data <= 8'b11111111;
		13'b0110110010101: data <= 8'b11111111;
		13'b0110110010110: data <= 8'b11111111;
		13'b0110110011001: data <= 8'b11111111;
		13'b0110110011010: data <= 8'b11111111;
		13'b0110110011011: data <= 8'b11111111;
		13'b0110110011100: data <= 8'b11111111;
		13'b0110110011101: data <= 8'b11111111;
		13'b0110111100001: data <= 8'b11111111;
		13'b0110111100010: data <= 8'b11111111;
		13'b0110111100011: data <= 8'b11111111;
		13'b0110111100100: data <= 8'b11111111;
		13'b0110111100101: data <= 8'b11111111;
		13'b0110111101010: data <= 8'b11111111;
		13'b0110111101011: data <= 8'b11111111;
		13'b0110111101100: data <= 8'b11111111;
		13'b0110111101101: data <= 8'b11111111;
		13'b0110111101110: data <= 8'b11111111;
		13'b0111000110000: data <= 8'b11111111;
		13'b0111000110001: data <= 8'b11111111;
		13'b0111000110010: data <= 8'b11111111;
		13'b0111000110011: data <= 8'b11111111;
		13'b0111000110100: data <= 8'b11111111;
		13'b0111000111011: data <= 8'b11111111;
		13'b0111000111100: data <= 8'b11111111;
		13'b0111000111101: data <= 8'b11111111;
		13'b0111000111110: data <= 8'b11111111;
		13'b0111000111111: data <= 8'b11111111;
		13'b0111001111111: data <= 8'b11111111;
		13'b0111010000000: data <= 8'b11111111;
		13'b0111010000001: data <= 8'b11111111;
		13'b0111010000010: data <= 8'b11111111;
		13'b0111010000011: data <= 8'b11111111;
		13'b0111010001100: data <= 8'b11111111;
		13'b0111010001101: data <= 8'b11111111;
		13'b0111010001110: data <= 8'b11111111;
		13'b0111010001111: data <= 8'b11111111;
		13'b0111010010000: data <= 8'b11111111;
		13'b0111011001110: data <= 8'b11111111;
		13'b0111011001111: data <= 8'b11111111;
		13'b0111011010000: data <= 8'b11111111;
		13'b0111011010001: data <= 8'b11111111;
		13'b0111011010010: data <= 8'b11111111;
		13'b0111011011101: data <= 8'b11111111;
		13'b0111011011110: data <= 8'b11111111;
		13'b0111011011111: data <= 8'b11111111;
		13'b0111011100000: data <= 8'b11111111;
		13'b0111011100001: data <= 8'b11111111;
		13'b0111100011101: data <= 8'b11111111;
		13'b0111100011110: data <= 8'b11111111;
		13'b0111100011111: data <= 8'b11111111;
		13'b0111100100000: data <= 8'b11111111;
		13'b0111100100001: data <= 8'b11111111;
		13'b0111100101110: data <= 8'b11111111;
		13'b0111100101111: data <= 8'b11111111;
		13'b0111100110000: data <= 8'b11111111;
		13'b0111100110001: data <= 8'b11111111;
		13'b0111100110010: data <= 8'b11111111;
		13'b0111101101100: data <= 8'b11111111;
		13'b0111101101101: data <= 8'b11111111;
		13'b0111101101110: data <= 8'b11111111;
		13'b0111101101111: data <= 8'b11111111;
		13'b0111101110000: data <= 8'b11111111;
		13'b0111101111111: data <= 8'b11111111;
		13'b0111110000000: data <= 8'b11111111;
		13'b0111110000001: data <= 8'b11111111;
		13'b0111110000010: data <= 8'b11111111;
		13'b0111110000011: data <= 8'b11111111;
		13'b0111110111011: data <= 8'b11111111;
		13'b0111110111100: data <= 8'b11111111;
		13'b0111110111101: data <= 8'b11111111;
		13'b0111110111110: data <= 8'b11111111;
		13'b0111110111111: data <= 8'b11111111;
		13'b0111111010000: data <= 8'b11111111;
		13'b0111111010001: data <= 8'b11111111;
		13'b0111111010010: data <= 8'b11111111;
		13'b0111111010011: data <= 8'b11111111;
		13'b0111111010100: data <= 8'b11111111;
		13'b1000000001010: data <= 8'b11111111;
		13'b1000000001011: data <= 8'b11111111;
		13'b1000000001100: data <= 8'b11111111;
		13'b1000000001101: data <= 8'b11111111;
		13'b1000000001110: data <= 8'b11111111;
		13'b1000000100001: data <= 8'b11111111;
		13'b1000000100010: data <= 8'b11111111;
		13'b1000000100011: data <= 8'b11111111;
		13'b1000000100100: data <= 8'b11111111;
		13'b1000000100101: data <= 8'b11111111;
		13'b1000001011001: data <= 8'b11111111;
		13'b1000001011010: data <= 8'b11111111;
		13'b1000001011011: data <= 8'b11111111;
		13'b1000001011100: data <= 8'b11111111;
		13'b1000001011101: data <= 8'b11111111;
		13'b1000001110010: data <= 8'b11111111;
		13'b1000001110011: data <= 8'b11111111;
		13'b1000001110100: data <= 8'b11111111;
		13'b1000001110101: data <= 8'b11111111;
		13'b1000001110110: data <= 8'b11111111;
		13'b1000010101000: data <= 8'b11111111;
		13'b1000010101001: data <= 8'b11111111;
		13'b1000010101010: data <= 8'b11111111;
		13'b1000010101011: data <= 8'b11111111;
		13'b1000010101100: data <= 8'b11111111;
		13'b1000011000011: data <= 8'b11111111;
		13'b1000011000100: data <= 8'b11111111;
		13'b1000011000101: data <= 8'b11111111;
		13'b1000011000110: data <= 8'b11111111;
		13'b1000011000111: data <= 8'b11111111;
		13'b1000011110111: data <= 8'b11111111;
		13'b1000011111000: data <= 8'b11111111;
		13'b1000011111001: data <= 8'b11111111;
		13'b1000011111010: data <= 8'b11111111;
		13'b1000011111011: data <= 8'b11111111;
		13'b1000100010100: data <= 8'b11111111;
		13'b1000100010101: data <= 8'b11111111;
		13'b1000100010110: data <= 8'b11111111;
		13'b1000100010111: data <= 8'b11111111;
		13'b1000100011000: data <= 8'b11111111;
		13'b1000101000110: data <= 8'b11111111;
		13'b1000101000111: data <= 8'b11111111;
		13'b1000101001000: data <= 8'b11111111;
		13'b1000101001001: data <= 8'b11111111;
		13'b1000101001010: data <= 8'b11111111;
		13'b1000101100101: data <= 8'b11111111;
		13'b1000101100110: data <= 8'b11111111;
		13'b1000101100111: data <= 8'b11111111;
		13'b1000101101000: data <= 8'b11111111;
		13'b1000101101001: data <= 8'b11111111;
		13'b1000110010101: data <= 8'b11111111;
		13'b1000110010110: data <= 8'b11111111;
		13'b1000110010111: data <= 8'b11111111;
		13'b1000110011000: data <= 8'b11111111;
		13'b1000110011001: data <= 8'b11111111;
		13'b1000110110110: data <= 8'b11111111;
		13'b1000110110111: data <= 8'b11111111;
		13'b1000110111000: data <= 8'b11111111;
		13'b1000110111001: data <= 8'b11111111;
		13'b1000110111010: data <= 8'b11111111;
		13'b1000111100100: data <= 8'b11111111;
		13'b1000111100101: data <= 8'b11111111;
		13'b1000111100110: data <= 8'b11111111;
		13'b1000111100111: data <= 8'b11111111;
		13'b1000111101000: data <= 8'b11111111;
		13'b1001000000111: data <= 8'b11111111;
		13'b1001000001000: data <= 8'b11111111;
		13'b1001000001001: data <= 8'b11111111;
		13'b1001000001010: data <= 8'b11111111;
		13'b1001000001011: data <= 8'b11111111;
		13'b1001000110011: data <= 8'b11111111;
		13'b1001000110100: data <= 8'b11111111;
		13'b1001000110101: data <= 8'b11111111;
		13'b1001000110110: data <= 8'b11111111;
		13'b1001000110111: data <= 8'b11111111;
		13'b1001001011000: data <= 8'b11111111;
		13'b1001001011001: data <= 8'b11111111;
		13'b1001001011010: data <= 8'b11111111;
		13'b1001001011011: data <= 8'b11111111;
		13'b1001001011100: data <= 8'b11111111;
		13'b1001010000010: data <= 8'b11111111;
		13'b1001010000011: data <= 8'b11111111;
		13'b1001010000100: data <= 8'b11111111;
		13'b1001010000101: data <= 8'b11111111;
		13'b1001010000110: data <= 8'b11111111;
		13'b1001010101001: data <= 8'b11111111;
		13'b1001010101010: data <= 8'b11111111;
		13'b1001010101011: data <= 8'b11111111;
		13'b1001010101100: data <= 8'b11111111;
		13'b1001010101101: data <= 8'b11111111;
		13'b1001011010001: data <= 8'b11111111;
		13'b1001011010010: data <= 8'b11111111;
		13'b1001011010011: data <= 8'b11111111;
		13'b1001011010100: data <= 8'b11111111;
		13'b1001011010101: data <= 8'b11111111;
		13'b1001011111010: data <= 8'b11111111;
		13'b1001011111011: data <= 8'b11111111;
		13'b1001011111100: data <= 8'b11111111;
		13'b1001011111101: data <= 8'b11111111;
		13'b1001011111110: data <= 8'b11111111;
		13'b1001100100000: data <= 8'b11111111;
		13'b1001100100001: data <= 8'b11111111;
		13'b1001100100010: data <= 8'b11111111;
		13'b1001100100011: data <= 8'b11111111;
		13'b1001100100100: data <= 8'b11111111;
		13'b1001101001011: data <= 8'b11111111;
		13'b1001101001100: data <= 8'b11111111;
		13'b1001101001101: data <= 8'b11111111;
		13'b1001101001110: data <= 8'b11111111;
		13'b1001101001111: data <= 8'b11111111;
		13'b1001101101111: data <= 8'b11111111;
		13'b1001101110000: data <= 8'b11111111;
		13'b1001101110001: data <= 8'b11111111;
		13'b1001101110010: data <= 8'b11111111;
		13'b1001101110011: data <= 8'b11111111;
		13'b1001110011100: data <= 8'b11111111;
		13'b1001110011101: data <= 8'b11111111;
		13'b1001110011110: data <= 8'b11111111;
		13'b1001110011111: data <= 8'b11111111;
		13'b1001110100000: data <= 8'b11111111;
		13'b1001110111110: data <= 8'b11111111;
		13'b1001110111111: data <= 8'b11111111;
		13'b1001111000000: data <= 8'b11111111;
		13'b1001111000001: data <= 8'b11111111;
		13'b1001111000010: data <= 8'b11111111;
		13'b1001111101101: data <= 8'b11111111;
		13'b1001111101110: data <= 8'b11111111;
		13'b1001111101111: data <= 8'b11111111;
		13'b1001111110000: data <= 8'b11111111;
		13'b1001111110001: data <= 8'b11111111;
		13'b1010000001110: data <= 8'b11111111;
		13'b1010000001111: data <= 8'b11111111;
		13'b1010000010000: data <= 8'b11111111;
		13'b1010000010001: data <= 8'b11111111;
		13'b1010000111110: data <= 8'b11111111;
		13'b1010000111111: data <= 8'b11111111;
		13'b1010001000000: data <= 8'b11111111;
		13'b1010001000001: data <= 8'b11111111;
		13'b1010001011111: data <= 8'b11111111;
		13'b1010001100000: data <= 8'b11111111;
		13'b1010010001111: data <= 8'b11111111;
		13'b1010010010000: data <= 8'b11111111;
		default: data <= 8'b00000000;
	endcase
end

endmodule
module digits_rom(
//inputs
clk, addr, 
//outputs
data);

(* rom_style = "block" *)

input wire clk;
input wire [7:0] addr;
output reg [7:0] data;

reg [7:0] addr_reg;

always @ (posedge clk)
	addr_reg <= addr;

always @ (*)
begin
	case(addr)
		8'b00000001: data <= 8'b11111111;
		8'b00000011: data <= 8'b11111111;
		8'b00000101: data <= 8'b11111111;
		8'b00000110: data <= 8'b11111111;
		8'b00001000: data <= 8'b11111111;
		8'b00001001: data <= 8'b11111111;
		8'b00001011: data <= 8'b11111111;
		8'b00001101: data <= 8'b11111111;
		8'b00010000: data <= 8'b11111111;
		8'b00010010: data <= 8'b11111111;
		8'b00010011: data <= 8'b11111111;
		8'b00010110: data <= 8'b11111111;
		8'b00011001: data <= 8'b11111111;
		8'b00011011: data <= 8'b11111111;
		8'b00011100: data <= 8'b11111111;
		8'b00011101: data <= 8'b11111111;
		8'b00011111: data <= 8'b11111111;
		8'b00100001: data <= 8'b11111111;
		8'b00100011: data <= 8'b11111111;
		8'b00100110: data <= 8'b11111111;
		8'b00101000: data <= 8'b11111111;
		8'b00101010: data <= 8'b11111111;
		8'b00101011: data <= 8'b11111111;
		8'b00101100: data <= 8'b11111111;
		8'b00101101: data <= 8'b11111111;
		8'b00101110: data <= 8'b11111111;
		8'b00110010: data <= 8'b11111111;
		8'b00110011: data <= 8'b11111111;
		8'b00110100: data <= 8'b11111111;
		8'b00111000: data <= 8'b11111111;
		8'b00111001: data <= 8'b11111111;
		8'b00111010: data <= 8'b11111111;
		8'b00111100: data <= 8'b11111111;
		8'b00111110: data <= 8'b11111111;
		8'b00111111: data <= 8'b11111111;
		8'b01000001: data <= 8'b11111111;
		8'b01000010: data <= 8'b11111111;
		8'b01000011: data <= 8'b11111111;
		8'b01000100: data <= 8'b11111111;
		8'b01000111: data <= 8'b11111111;
		8'b01001010: data <= 8'b11111111;
		8'b01001011: data <= 8'b11111111;
		8'b01001100: data <= 8'b11111111;
		8'b01001101: data <= 8'b11111111;
		8'b01001110: data <= 8'b11111111;
		8'b01010001: data <= 8'b11111111;
		8'b01010010: data <= 8'b11111111;
		8'b01010110: data <= 8'b11111111;
		8'b01010111: data <= 8'b11111111;
		8'b01011000: data <= 8'b11111111;
		8'b01011011: data <= 8'b11111111;
		8'b01011100: data <= 8'b11111111;
		8'b01011101: data <= 8'b11111111;
		8'b01100000: data <= 8'b11111111;
		8'b01100001: data <= 8'b11111111;
		8'b01100011: data <= 8'b11111111;
		8'b01100101: data <= 8'b11111111;
		8'b01100111: data <= 8'b11111111;
		8'b01101001: data <= 8'b11111111;
		8'b01101010: data <= 8'b11111111;
		8'b01101011: data <= 8'b11111111;
		8'b01101110: data <= 8'b11111111;
		8'b01110000: data <= 8'b11111111;
		8'b01110010: data <= 8'b11111111;
		8'b01110101: data <= 8'b11111111;
		8'b01111001: data <= 8'b11111111;
		8'b01111011: data <= 8'b11111111;
		8'b01111101: data <= 8'b11111111;
		8'b01111111: data <= 8'b11111111;
		8'b10000001: data <= 8'b11111111;
		8'b10000011: data <= 8'b11111111;
		8'b10000101: data <= 8'b11111111;
		8'b10001000: data <= 8'b11111111;
		8'b10001010: data <= 8'b11111111;
		8'b10001100: data <= 8'b11111111;
		8'b10001110: data <= 8'b11111111;
		8'b10001111: data <= 8'b11111111;
		8'b10010010: data <= 8'b11111111;
		8'b10010101: data <= 8'b11111111;
		default: data <= 8'b00000000;
	endcase
end

endmodule